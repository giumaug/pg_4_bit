magic
tech sky130A
timestamp 1738578133
<< metal1 >>
rect 100 20245 925 20255
rect 100 20205 110 20245
rect 150 20205 170 20245
rect 210 20205 230 20245
rect 270 20205 925 20245
rect 100 20195 925 20205
rect 400 19975 925 19985
rect 400 19935 410 19975
rect 450 19935 470 19975
rect 510 19935 530 19975
rect 570 19935 925 19975
rect 400 19925 925 19935
<< via1 >>
rect 110 20205 150 20245
rect 170 20205 210 20245
rect 230 20205 270 20245
rect 410 19935 450 19975
rect 470 19935 510 19975
rect 530 19935 570 19975
<< metal2 >>
rect 100 20245 300 20255
rect 100 20205 110 20245
rect 150 20205 170 20245
rect 210 20205 230 20245
rect 270 20205 300 20245
rect 100 20195 300 20205
rect 400 19975 600 19985
rect 400 19935 410 19975
rect 450 19935 470 19975
rect 510 19935 530 19975
rect 570 19935 600 19975
rect 400 19925 600 19935
<< via2 >>
rect 110 20205 150 20245
rect 170 20205 210 20245
rect 230 20205 270 20245
rect 410 19935 450 19975
rect 470 19935 510 19975
rect 530 19935 570 19975
<< metal3 >>
rect 400 21990 945 22000
rect 400 21950 410 21990
rect 450 21950 470 21990
rect 510 21950 530 21990
rect 570 21951 945 21990
rect 570 21950 600 21951
rect 815 21950 945 21951
rect 400 21935 600 21950
rect 100 20245 300 20255
rect 100 20205 110 20245
rect 150 20205 170 20245
rect 210 20205 230 20245
rect 270 20205 300 20245
rect 100 20195 300 20205
rect 400 19975 600 19985
rect 400 19935 410 19975
rect 450 19935 470 19975
rect 510 19935 530 19975
rect 570 19935 600 19975
rect 400 19925 600 19935
<< via3 >>
rect 410 21950 450 21990
rect 470 21950 510 21990
rect 530 21950 570 21990
rect 110 20205 150 20245
rect 170 20205 210 20245
rect 230 20205 270 20245
rect 410 19935 450 19975
rect 470 19935 510 19975
rect 530 19935 570 19975
<< metal4 >>
rect 3067 22490 3097 22576
rect 3343 22495 3373 22576
rect 3619 22495 3649 22576
rect 3895 22495 3925 22576
rect 4171 22495 4201 22576
rect 100 20245 300 22076
rect 100 20205 110 20245
rect 150 20205 170 20245
rect 210 20205 230 20245
rect 270 20205 300 20245
rect 100 500 300 20205
rect 400 21990 600 22076
rect 3060 22030 3105 22490
rect 3340 22035 3385 22495
rect 3615 22035 3660 22495
rect 3890 21990 3935 22495
rect 4170 21990 4210 22495
rect 4447 22490 4477 22576
rect 4445 22000 4485 22490
rect 4723 22485 4753 22576
rect 4999 22490 5029 22576
rect 4720 21995 4760 22485
rect 4995 22000 5035 22490
rect 5275 22485 5305 22576
rect 5551 22490 5581 22576
rect 5827 22490 5857 22576
rect 5270 21995 5310 22485
rect 5550 22000 5590 22490
rect 5825 22000 5865 22490
rect 6103 22485 6133 22576
rect 6379 22490 6409 22576
rect 6655 22490 6685 22576
rect 6931 22490 6961 22576
rect 7207 22490 7237 22576
rect 7483 22490 7513 22576
rect 7759 22490 7789 22576
rect 8035 22490 8065 22576
rect 8311 22490 8341 22576
rect 8587 22490 8617 22576
rect 8863 22490 8893 22576
rect 9139 22495 9169 22576
rect 9415 22495 9445 22576
rect 6100 21995 6140 22485
rect 6375 22000 6415 22490
rect 6650 22000 6690 22490
rect 6930 22000 6970 22490
rect 7205 22000 7245 22490
rect 7480 22040 7520 22490
rect 7755 22035 7795 22490
rect 8030 22035 8070 22490
rect 8310 22035 8350 22490
rect 8580 22030 8625 22490
rect 8860 22030 8905 22490
rect 9130 22030 9175 22495
rect 9410 22030 9455 22495
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22490 11929 22576
rect 12175 22490 12205 22576
rect 12451 22570 12481 22576
rect 11895 22035 11940 22490
rect 400 21950 410 21990
rect 450 21950 470 21990
rect 510 21950 530 21990
rect 570 21950 600 21990
rect 400 19975 600 21950
rect 12175 21820 12215 22490
rect 12450 21900 12490 22570
rect 12727 22490 12757 22576
rect 13003 22490 13033 22576
rect 13279 22490 13309 22576
rect 13555 22490 13585 22576
rect 13831 22490 13861 22576
rect 12725 22030 12770 22490
rect 13000 22030 13045 22490
rect 13270 22030 13315 22490
rect 13550 22030 13595 22490
rect 13820 22030 13865 22490
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 400 19935 410 19975
rect 450 19935 470 19975
rect 510 19935 530 19975
rect 570 19935 600 19975
rect 400 500 600 19935
use cell  cell_0
timestamp 1738491202
transform 1 0 3 0 1 11080
box 908 8845 14700 10967
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 100 500 300 22076 1 FreeSans 2 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 2 0 0 0 VGND
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
