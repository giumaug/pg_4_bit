VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_pg_4_bit
  CLASS BLOCK ;
  FOREIGN tt_um_pg_4_bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 110.520 144.130 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 110.520 146.890 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 110.520 141.370 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 101.600 147.000 102.100 ;
      LAYER via3 ;
        RECT 138.200 101.650 138.600 102.050 ;
      LAYER met4 ;
        RECT 138.310 110.850 138.610 111.520 ;
        RECT 138.200 110.520 138.610 110.850 ;
        RECT 138.200 102.100 138.600 110.520 ;
        RECT 138.100 101.600 138.650 102.100 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 102.500 147.000 103.000 ;
      LAYER via3 ;
        RECT 135.500 102.550 135.900 102.950 ;
      LAYER met4 ;
        RECT 135.550 110.600 135.850 111.520 ;
        RECT 135.500 103.000 135.900 110.600 ;
        RECT 135.400 102.500 135.950 103.000 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 103.400 147.000 103.900 ;
      LAYER via3 ;
        RECT 132.700 103.450 133.100 103.850 ;
      LAYER met4 ;
        RECT 132.790 110.600 133.090 111.520 ;
        RECT 132.700 103.900 133.100 110.600 ;
        RECT 132.600 103.400 133.150 103.900 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 104.300 147.000 104.800 ;
      LAYER via3 ;
        RECT 130.000 104.350 130.400 104.750 ;
      LAYER met4 ;
        RECT 130.030 110.600 130.330 111.520 ;
        RECT 130.000 104.800 130.400 110.600 ;
        RECT 129.900 104.300 130.450 104.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 105.200 147.000 105.700 ;
      LAYER via3 ;
        RECT 127.250 105.240 127.650 105.650 ;
      LAYER met4 ;
        RECT 127.270 110.650 127.570 111.520 ;
        RECT 127.250 105.700 127.650 110.650 ;
        RECT 127.150 105.200 127.700 105.700 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 124.400 106.500 124.950 106.550 ;
        RECT 80.500 106.100 147.000 106.500 ;
        RECT 124.400 106.050 124.950 106.100 ;
      LAYER via3 ;
        RECT 124.400 106.100 124.900 106.500 ;
      LAYER met4 ;
        RECT 124.510 110.600 124.810 111.520 ;
        RECT 124.500 106.550 124.850 110.600 ;
        RECT 124.350 106.050 124.950 106.550 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 106.900 147.000 107.400 ;
      LAYER via3 ;
        RECT 121.700 106.950 122.050 107.350 ;
      LAYER met4 ;
        RECT 121.750 107.400 122.050 111.520 ;
        RECT 121.650 106.900 122.100 107.400 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 107.800 147.000 108.300 ;
      LAYER via3 ;
        RECT 118.900 107.850 119.300 108.250 ;
      LAYER met4 ;
        RECT 118.990 110.600 119.290 111.520 ;
        RECT 118.950 108.300 119.300 110.600 ;
        RECT 118.850 107.800 119.350 108.300 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 110.520 116.530 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 110.520 113.770 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 110.520 111.010 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 110.520 108.250 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 110.520 105.490 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 110.520 102.730 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 110.520 99.970 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 110.520 97.210 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met3 ;
        RECT 80.500 108.700 147.000 109.200 ;
      LAYER met4 ;
        RECT 4.000 112.880 6.000 220.760 ;
        RECT 49.990 110.520 50.290 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 47.230 110.520 47.530 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 44.470 110.520 44.770 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 41.710 110.520 42.010 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 38.950 110.520 39.250 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 36.190 110.520 36.490 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 33.430 110.520 33.730 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 30.670 110.520 30.970 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 72.070 110.520 72.370 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 69.310 110.520 69.610 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 66.550 110.520 66.850 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 63.790 110.520 64.090 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 61.030 110.520 61.330 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 58.270 110.520 58.570 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 55.510 110.520 55.810 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.193650 ;
    PORT
      LAYER met4 ;
        RECT 52.750 110.520 53.050 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.657000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 94.400 147.000 94.900 ;
      LAYER via3 ;
        RECT 94.100 94.450 94.500 94.850 ;
      LAYER met4 ;
        RECT 94.150 110.600 94.450 111.520 ;
        RECT 94.100 94.900 94.500 110.600 ;
        RECT 94.050 94.400 94.550 94.900 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met3 ;
        RECT 80.500 95.300 147.000 95.800 ;
      LAYER via3 ;
        RECT 91.300 95.350 91.700 95.750 ;
      LAYER met4 ;
        RECT 91.390 110.600 91.690 111.520 ;
        RECT 91.300 95.800 91.700 110.600 ;
        RECT 91.250 95.300 91.750 95.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.657000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 96.200 147.000 96.700 ;
      LAYER via3 ;
        RECT 88.600 96.250 89.000 96.650 ;
      LAYER met4 ;
        RECT 88.630 110.600 88.930 111.520 ;
        RECT 88.600 96.700 89.000 110.600 ;
        RECT 88.550 96.200 89.050 96.700 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met3 ;
        RECT 80.500 97.100 147.000 97.600 ;
      LAYER via3 ;
        RECT 85.800 97.150 86.200 97.550 ;
      LAYER met4 ;
        RECT 85.870 110.600 86.170 111.520 ;
        RECT 85.800 97.600 86.200 110.600 ;
        RECT 85.750 97.100 86.250 97.600 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.657000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 98.000 147.000 98.500 ;
      LAYER via3 ;
        RECT 83.100 98.050 83.450 98.450 ;
      LAYER met4 ;
        RECT 83.110 110.600 83.410 111.520 ;
        RECT 83.100 98.500 83.450 110.600 ;
        RECT 83.050 98.000 83.500 98.500 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met3 ;
        RECT 80.500 98.900 147.000 99.400 ;
      LAYER via3 ;
        RECT 80.500 98.950 80.650 99.350 ;
      LAYER met4 ;
        RECT 80.350 110.520 80.650 111.520 ;
        RECT 80.500 99.400 80.650 110.520 ;
        RECT 80.500 98.900 80.700 99.400 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.657000 ;
    PORT
      LAYER met3 ;
        RECT 80.500 99.800 147.000 100.300 ;
      LAYER met4 ;
        RECT 77.590 110.520 77.890 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met3 ;
        RECT 80.500 100.700 147.000 101.200 ;
      LAYER met4 ;
        RECT 74.830 110.520 75.130 111.520 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 34.400 90.045 60.740 91.650 ;
      LAYER pwell ;
        RECT 35.735 89.750 36.685 89.755 ;
        RECT 37.385 89.750 40.555 89.755 ;
        RECT 35.735 89.665 40.555 89.750 ;
        RECT 42.135 89.750 43.085 89.755 ;
        RECT 43.785 89.750 46.955 89.755 ;
        RECT 42.135 89.715 46.955 89.750 ;
        RECT 49.325 89.750 50.275 89.755 ;
        RECT 50.975 89.750 54.145 89.755 ;
        RECT 42.135 89.665 47.785 89.715 ;
        RECT 49.325 89.665 54.145 89.750 ;
        RECT 55.725 89.665 60.545 89.755 ;
        RECT 34.755 88.980 60.545 89.665 ;
        RECT 34.755 88.975 43.085 88.980 ;
        RECT 34.755 88.845 36.685 88.975 ;
        RECT 37.385 88.845 40.555 88.975 ;
        RECT 41.155 88.845 43.085 88.975 ;
        RECT 43.785 88.975 47.785 88.980 ;
        RECT 43.785 88.845 46.955 88.975 ;
        RECT 47.355 88.930 47.785 88.975 ;
        RECT 48.345 88.975 54.145 88.980 ;
        RECT 48.345 88.845 50.275 88.975 ;
        RECT 50.975 88.845 54.145 88.975 ;
        RECT 54.745 88.845 56.675 88.980 ;
        RECT 57.375 88.845 60.545 88.980 ;
        RECT 34.755 88.825 34.905 88.845 ;
        RECT 34.735 88.655 34.905 88.825 ;
        RECT 37.485 88.655 37.655 88.845 ;
        RECT 41.155 88.825 41.305 88.845 ;
        RECT 41.135 88.655 41.305 88.825 ;
        RECT 43.885 88.655 44.055 88.845 ;
        RECT 48.345 88.825 48.495 88.845 ;
        RECT 48.325 88.655 48.495 88.825 ;
        RECT 51.075 88.655 51.245 88.845 ;
        RECT 54.745 88.825 54.895 88.845 ;
        RECT 54.725 88.655 54.895 88.825 ;
        RECT 57.475 88.655 57.645 88.845 ;
      LAYER li1 ;
        RECT 34.590 91.375 60.550 91.545 ;
        RECT 34.875 90.705 35.155 91.375 ;
        RECT 35.325 90.485 35.625 91.035 ;
        RECT 35.825 90.655 36.155 91.375 ;
        RECT 36.345 90.655 36.805 91.205 ;
        RECT 34.690 90.065 34.955 90.425 ;
        RECT 35.325 90.315 36.265 90.485 ;
        RECT 36.095 90.065 36.265 90.315 ;
        RECT 34.690 89.815 35.365 90.065 ;
        RECT 35.585 89.815 35.925 90.065 ;
        RECT 36.095 89.735 36.385 90.065 ;
        RECT 36.095 89.645 36.265 89.735 ;
        RECT 34.875 89.455 36.265 89.645 ;
        RECT 34.875 89.095 35.205 89.455 ;
        RECT 36.555 89.285 36.805 90.655 ;
        RECT 37.425 90.525 37.805 91.205 ;
        RECT 38.395 90.525 38.565 91.375 ;
        RECT 38.735 90.695 39.065 91.205 ;
        RECT 39.235 90.865 39.405 91.375 ;
        RECT 39.575 90.695 39.975 91.205 ;
        RECT 38.735 90.525 39.975 90.695 ;
        RECT 37.425 89.565 37.595 90.525 ;
        RECT 37.765 90.185 39.070 90.355 ;
        RECT 40.155 90.275 40.475 91.205 ;
        RECT 41.275 90.705 41.555 91.375 ;
        RECT 41.725 90.485 42.025 91.035 ;
        RECT 42.225 90.655 42.555 91.375 ;
        RECT 42.745 90.655 43.205 91.205 ;
        RECT 37.765 89.735 38.010 90.185 ;
        RECT 38.180 89.815 38.730 90.015 ;
        RECT 38.900 89.985 39.070 90.185 ;
        RECT 39.845 90.105 40.475 90.275 ;
        RECT 38.900 89.815 39.275 89.985 ;
        RECT 39.445 89.565 39.675 90.065 ;
        RECT 37.425 89.395 39.675 89.565 ;
        RECT 35.825 88.825 36.075 89.285 ;
        RECT 36.245 88.995 36.805 89.285 ;
        RECT 37.475 88.825 37.805 89.215 ;
        RECT 37.975 89.075 38.145 89.395 ;
        RECT 39.845 89.225 40.015 90.105 ;
        RECT 41.090 90.065 41.355 90.425 ;
        RECT 41.725 90.315 42.665 90.485 ;
        RECT 42.495 90.065 42.665 90.315 ;
        RECT 41.090 89.815 41.765 90.065 ;
        RECT 41.985 89.815 42.325 90.065 ;
        RECT 42.495 89.735 42.785 90.065 ;
        RECT 38.315 88.825 38.645 89.215 ;
        RECT 39.060 89.055 40.015 89.225 ;
        RECT 40.185 88.825 40.475 89.660 ;
        RECT 42.495 89.645 42.665 89.735 ;
        RECT 41.275 89.455 42.665 89.645 ;
        RECT 41.275 89.095 41.605 89.455 ;
        RECT 42.955 89.285 43.205 90.655 ;
        RECT 43.825 90.525 44.205 91.205 ;
        RECT 44.795 90.525 44.965 91.375 ;
        RECT 45.135 90.695 45.465 91.205 ;
        RECT 45.635 90.865 45.805 91.375 ;
        RECT 45.975 90.695 46.375 91.205 ;
        RECT 45.135 90.525 46.375 90.695 ;
        RECT 43.825 89.565 43.995 90.525 ;
        RECT 44.165 90.185 45.470 90.355 ;
        RECT 46.555 90.275 46.875 91.205 ;
        RECT 44.165 89.735 44.410 90.185 ;
        RECT 44.580 89.815 45.130 90.015 ;
        RECT 45.300 89.985 45.470 90.185 ;
        RECT 46.245 90.105 46.875 90.275 ;
        RECT 47.425 90.210 47.715 91.375 ;
        RECT 48.465 90.705 48.745 91.375 ;
        RECT 48.915 90.485 49.215 91.035 ;
        RECT 49.415 90.655 49.745 91.375 ;
        RECT 49.935 90.655 50.395 91.205 ;
        RECT 45.300 89.815 45.675 89.985 ;
        RECT 45.845 89.565 46.075 90.065 ;
        RECT 43.825 89.395 46.075 89.565 ;
        RECT 42.225 88.825 42.475 89.285 ;
        RECT 42.645 88.995 43.205 89.285 ;
        RECT 43.875 88.825 44.205 89.215 ;
        RECT 44.375 89.075 44.545 89.395 ;
        RECT 46.245 89.225 46.415 90.105 ;
        RECT 48.280 90.065 48.545 90.425 ;
        RECT 48.915 90.315 49.855 90.485 ;
        RECT 49.685 90.065 49.855 90.315 ;
        RECT 48.280 89.815 48.955 90.065 ;
        RECT 49.175 89.815 49.515 90.065 ;
        RECT 49.685 89.735 49.975 90.065 ;
        RECT 44.715 88.825 45.045 89.215 ;
        RECT 45.460 89.055 46.415 89.225 ;
        RECT 46.585 88.825 46.875 89.660 ;
        RECT 49.685 89.645 49.855 89.735 ;
        RECT 47.425 88.825 47.715 89.550 ;
        RECT 48.465 89.455 49.855 89.645 ;
        RECT 48.465 89.095 48.795 89.455 ;
        RECT 50.145 89.285 50.395 90.655 ;
        RECT 51.015 90.525 51.395 91.205 ;
        RECT 51.985 90.525 52.155 91.375 ;
        RECT 52.325 90.695 52.655 91.205 ;
        RECT 52.825 90.865 52.995 91.375 ;
        RECT 53.165 90.695 53.565 91.205 ;
        RECT 52.325 90.525 53.565 90.695 ;
        RECT 51.015 89.565 51.185 90.525 ;
        RECT 51.355 90.185 52.660 90.355 ;
        RECT 53.745 90.275 54.065 91.205 ;
        RECT 54.865 90.705 55.145 91.375 ;
        RECT 55.315 90.485 55.615 91.035 ;
        RECT 55.815 90.655 56.145 91.375 ;
        RECT 56.335 90.655 56.795 91.205 ;
        RECT 51.355 89.735 51.600 90.185 ;
        RECT 51.770 89.815 52.320 90.015 ;
        RECT 52.490 89.985 52.660 90.185 ;
        RECT 53.435 90.105 54.065 90.275 ;
        RECT 52.490 89.815 52.865 89.985 ;
        RECT 53.035 89.565 53.265 90.065 ;
        RECT 51.015 89.395 53.265 89.565 ;
        RECT 49.415 88.825 49.665 89.285 ;
        RECT 49.835 88.995 50.395 89.285 ;
        RECT 51.065 88.825 51.395 89.215 ;
        RECT 51.565 89.075 51.735 89.395 ;
        RECT 53.435 89.225 53.605 90.105 ;
        RECT 54.680 90.065 54.945 90.425 ;
        RECT 55.315 90.315 56.255 90.485 ;
        RECT 56.085 90.065 56.255 90.315 ;
        RECT 54.680 89.815 55.355 90.065 ;
        RECT 55.575 89.815 55.915 90.065 ;
        RECT 56.085 89.735 56.375 90.065 ;
        RECT 51.905 88.825 52.235 89.215 ;
        RECT 52.650 89.055 53.605 89.225 ;
        RECT 53.775 88.825 54.065 89.660 ;
        RECT 56.085 89.645 56.255 89.735 ;
        RECT 54.865 89.455 56.255 89.645 ;
        RECT 54.865 89.095 55.195 89.455 ;
        RECT 56.545 89.285 56.795 90.655 ;
        RECT 57.415 90.525 57.795 91.205 ;
        RECT 58.385 90.525 58.555 91.375 ;
        RECT 58.725 90.695 59.055 91.205 ;
        RECT 59.225 90.865 59.395 91.375 ;
        RECT 59.565 90.695 59.965 91.205 ;
        RECT 58.725 90.525 59.965 90.695 ;
        RECT 57.415 89.565 57.585 90.525 ;
        RECT 57.755 90.185 59.060 90.355 ;
        RECT 60.145 90.275 60.465 91.205 ;
        RECT 57.755 89.735 58.000 90.185 ;
        RECT 58.170 89.815 58.720 90.015 ;
        RECT 58.890 89.985 59.060 90.185 ;
        RECT 59.835 90.105 60.465 90.275 ;
        RECT 58.890 89.815 59.265 89.985 ;
        RECT 59.435 89.565 59.665 90.065 ;
        RECT 57.415 89.395 59.665 89.565 ;
        RECT 55.815 88.825 56.065 89.285 ;
        RECT 56.235 88.995 56.795 89.285 ;
        RECT 57.465 88.825 57.795 89.215 ;
        RECT 57.965 89.075 58.135 89.395 ;
        RECT 59.835 89.225 60.005 90.105 ;
        RECT 58.305 88.825 58.635 89.215 ;
        RECT 59.050 89.055 60.005 89.225 ;
        RECT 60.175 88.825 60.465 89.660 ;
        RECT 34.590 88.655 60.550 88.825 ;
        RECT 36.785 88.650 37.375 88.655 ;
      LAYER mcon ;
        RECT 34.735 91.375 34.905 91.545 ;
        RECT 35.195 91.375 35.365 91.545 ;
        RECT 35.655 91.375 35.825 91.545 ;
        RECT 36.115 91.375 36.285 91.545 ;
        RECT 36.575 91.375 36.745 91.545 ;
        RECT 37.020 91.375 37.200 91.545 ;
        RECT 37.485 91.375 37.655 91.545 ;
        RECT 37.945 91.375 38.115 91.545 ;
        RECT 38.405 91.375 38.575 91.545 ;
        RECT 38.865 91.375 39.035 91.545 ;
        RECT 39.325 91.375 39.495 91.545 ;
        RECT 39.785 91.375 39.955 91.545 ;
        RECT 40.245 91.375 40.415 91.545 ;
        RECT 40.700 91.375 40.875 91.545 ;
        RECT 41.135 91.375 41.305 91.545 ;
        RECT 41.595 91.375 41.765 91.545 ;
        RECT 42.055 91.375 42.225 91.545 ;
        RECT 42.515 91.375 42.685 91.545 ;
        RECT 42.975 91.375 43.145 91.545 ;
        RECT 43.420 91.375 43.600 91.545 ;
        RECT 43.885 91.375 44.055 91.545 ;
        RECT 44.345 91.375 44.515 91.545 ;
        RECT 44.805 91.375 44.975 91.545 ;
        RECT 45.265 91.375 45.435 91.545 ;
        RECT 45.725 91.375 45.895 91.545 ;
        RECT 46.185 91.375 46.355 91.545 ;
        RECT 46.645 91.375 46.815 91.545 ;
        RECT 47.050 91.375 47.225 91.545 ;
        RECT 47.485 91.375 47.655 91.545 ;
        RECT 47.925 91.375 48.100 91.545 ;
        RECT 48.325 91.375 48.495 91.545 ;
        RECT 48.785 91.375 48.955 91.545 ;
        RECT 49.245 91.375 49.415 91.545 ;
        RECT 49.705 91.375 49.875 91.545 ;
        RECT 50.165 91.375 50.335 91.545 ;
        RECT 50.615 91.375 50.790 91.545 ;
        RECT 51.075 91.375 51.245 91.545 ;
        RECT 51.535 91.375 51.705 91.545 ;
        RECT 51.995 91.375 52.165 91.545 ;
        RECT 52.455 91.375 52.625 91.545 ;
        RECT 52.915 91.375 53.085 91.545 ;
        RECT 53.375 91.375 53.545 91.545 ;
        RECT 53.835 91.375 54.005 91.545 ;
        RECT 54.290 91.375 54.465 91.545 ;
        RECT 54.725 91.375 54.895 91.545 ;
        RECT 55.185 91.375 55.355 91.545 ;
        RECT 55.645 91.375 55.815 91.545 ;
        RECT 56.105 91.375 56.275 91.545 ;
        RECT 56.565 91.375 56.735 91.545 ;
        RECT 57.015 91.375 57.190 91.545 ;
        RECT 57.475 91.375 57.645 91.545 ;
        RECT 57.935 91.375 58.105 91.545 ;
        RECT 58.395 91.375 58.565 91.545 ;
        RECT 58.855 91.375 59.025 91.545 ;
        RECT 59.315 91.375 59.485 91.545 ;
        RECT 59.775 91.375 59.945 91.545 ;
        RECT 60.235 91.375 60.405 91.545 ;
        RECT 36.425 90.655 36.595 90.825 ;
        RECT 34.960 89.815 35.130 89.985 ;
        RECT 35.665 89.815 35.835 89.985 ;
        RECT 40.175 90.275 40.345 90.445 ;
        RECT 42.825 90.655 42.995 90.825 ;
        RECT 37.765 89.815 37.935 89.985 ;
        RECT 38.350 89.815 38.520 89.985 ;
        RECT 41.360 89.815 41.530 89.985 ;
        RECT 42.065 89.815 42.235 89.985 ;
        RECT 46.575 90.615 46.745 90.785 ;
        RECT 44.165 89.815 44.335 89.985 ;
        RECT 44.750 89.815 44.920 89.985 ;
        RECT 50.015 90.655 50.185 90.825 ;
        RECT 48.550 89.815 48.720 89.985 ;
        RECT 49.255 89.815 49.425 89.985 ;
        RECT 53.765 90.275 53.935 90.445 ;
        RECT 56.415 90.655 56.585 90.825 ;
        RECT 51.940 89.815 52.110 89.985 ;
        RECT 52.615 89.815 52.785 89.985 ;
        RECT 54.950 89.815 55.120 89.985 ;
        RECT 55.655 89.815 55.825 89.985 ;
        RECT 60.165 90.615 60.335 90.785 ;
        RECT 57.755 89.815 57.925 89.985 ;
        RECT 58.340 89.815 58.510 89.985 ;
        RECT 34.735 88.655 34.905 88.825 ;
        RECT 35.195 88.655 35.365 88.825 ;
        RECT 35.655 88.655 35.825 88.825 ;
        RECT 36.115 88.655 36.285 88.825 ;
        RECT 36.575 88.655 36.745 88.825 ;
        RECT 37.020 88.650 37.200 88.825 ;
        RECT 37.485 88.655 37.655 88.825 ;
        RECT 37.945 88.655 38.115 88.825 ;
        RECT 38.405 88.655 38.575 88.825 ;
        RECT 38.865 88.655 39.035 88.825 ;
        RECT 39.325 88.655 39.495 88.825 ;
        RECT 39.785 88.655 39.955 88.825 ;
        RECT 40.245 88.655 40.415 88.825 ;
        RECT 40.670 88.655 40.850 88.825 ;
        RECT 41.135 88.655 41.305 88.825 ;
        RECT 41.595 88.655 41.765 88.825 ;
        RECT 42.055 88.655 42.225 88.825 ;
        RECT 42.515 88.655 42.685 88.825 ;
        RECT 42.975 88.655 43.145 88.825 ;
        RECT 43.425 88.655 43.600 88.825 ;
        RECT 43.885 88.655 44.055 88.825 ;
        RECT 44.345 88.655 44.515 88.825 ;
        RECT 44.805 88.655 44.975 88.825 ;
        RECT 45.265 88.655 45.435 88.825 ;
        RECT 45.725 88.655 45.895 88.825 ;
        RECT 46.185 88.655 46.355 88.825 ;
        RECT 46.645 88.655 46.815 88.825 ;
        RECT 47.050 88.655 47.225 88.825 ;
        RECT 47.485 88.655 47.655 88.825 ;
        RECT 47.900 88.655 48.075 88.825 ;
        RECT 48.325 88.655 48.495 88.825 ;
        RECT 48.785 88.655 48.955 88.825 ;
        RECT 49.245 88.655 49.415 88.825 ;
        RECT 49.705 88.655 49.875 88.825 ;
        RECT 50.165 88.655 50.335 88.825 ;
        RECT 50.615 88.655 50.790 88.825 ;
        RECT 51.075 88.655 51.245 88.825 ;
        RECT 51.535 88.655 51.705 88.825 ;
        RECT 51.995 88.655 52.165 88.825 ;
        RECT 52.455 88.655 52.625 88.825 ;
        RECT 52.915 88.655 53.085 88.825 ;
        RECT 53.375 88.655 53.545 88.825 ;
        RECT 53.835 88.655 54.005 88.825 ;
        RECT 54.290 88.655 54.465 88.825 ;
        RECT 54.725 88.655 54.895 88.825 ;
        RECT 55.185 88.655 55.355 88.825 ;
        RECT 55.645 88.655 55.815 88.825 ;
        RECT 56.105 88.655 56.275 88.825 ;
        RECT 56.565 88.655 56.735 88.825 ;
        RECT 57.015 88.655 57.190 88.825 ;
        RECT 57.475 88.655 57.645 88.825 ;
        RECT 57.935 88.655 58.105 88.825 ;
        RECT 58.395 88.655 58.565 88.825 ;
        RECT 58.855 88.655 59.025 88.825 ;
        RECT 59.315 88.655 59.485 88.825 ;
        RECT 59.775 88.655 59.945 88.825 ;
        RECT 60.235 88.655 60.405 88.825 ;
      LAYER met1 ;
        RECT 1.000 91.700 34.700 91.750 ;
        RECT 1.000 91.220 60.550 91.700 ;
        RECT 1.000 91.175 34.700 91.220 ;
        RECT 36.300 90.875 36.750 91.000 ;
        RECT 42.700 90.875 43.150 91.000 ;
        RECT 36.300 90.625 36.800 90.875 ;
        RECT 42.700 90.625 43.200 90.875 ;
        RECT 36.300 90.550 36.750 90.625 ;
        RECT 34.900 90.255 38.600 90.400 ;
        RECT 34.900 90.250 37.970 90.255 ;
        RECT 34.900 90.150 35.250 90.250 ;
        RECT 34.800 89.700 35.250 90.150 ;
        RECT 35.600 89.800 35.900 90.050 ;
        RECT 35.585 89.700 35.900 89.800 ;
        RECT 37.650 89.700 38.100 90.100 ;
        RECT 38.250 89.750 38.600 90.255 ;
        RECT 40.100 90.150 40.550 90.600 ;
        RECT 42.700 90.550 43.150 90.625 ;
        RECT 46.450 90.500 46.950 90.950 ;
        RECT 49.900 90.875 50.350 91.000 ;
        RECT 56.300 90.875 56.750 91.000 ;
        RECT 49.900 90.595 50.365 90.875 ;
        RECT 56.300 90.600 56.790 90.875 ;
        RECT 49.900 90.550 50.350 90.595 ;
        RECT 41.300 90.250 45.000 90.400 ;
        RECT 41.300 90.100 41.600 90.250 ;
        RECT 35.585 89.650 38.100 89.700 ;
        RECT 41.200 89.650 41.650 90.100 ;
        RECT 42.000 89.750 42.300 90.050 ;
        RECT 35.585 89.550 38.000 89.650 ;
        RECT 42.000 89.600 42.150 89.750 ;
        RECT 44.050 89.600 44.500 90.100 ;
        RECT 44.700 89.750 45.000 90.250 ;
        RECT 48.490 90.250 52.140 90.400 ;
        RECT 48.490 90.100 48.790 90.250 ;
        RECT 48.400 89.650 48.850 90.100 ;
        RECT 42.000 89.455 44.500 89.600 ;
        RECT 42.300 89.450 44.500 89.455 ;
        RECT 49.190 89.600 49.490 90.050 ;
        RECT 51.890 89.750 52.140 90.250 ;
        RECT 53.650 90.150 54.100 90.600 ;
        RECT 56.300 90.550 56.750 90.600 ;
        RECT 60.050 90.450 60.500 90.900 ;
        RECT 54.890 90.250 58.590 90.400 ;
        RECT 52.450 89.700 52.900 90.150 ;
        RECT 54.890 90.100 55.190 90.250 ;
        RECT 52.450 89.600 52.840 89.700 ;
        RECT 54.800 89.650 55.250 90.100 ;
        RECT 49.190 89.450 52.840 89.600 ;
        RECT 55.590 89.600 55.890 90.050 ;
        RECT 57.600 89.600 58.050 90.100 ;
        RECT 58.290 89.750 58.590 90.250 ;
        RECT 55.590 89.450 58.050 89.600 ;
        RECT 4.000 88.980 34.675 89.025 ;
        RECT 4.000 88.975 36.890 88.980 ;
        RECT 37.340 88.975 60.550 88.980 ;
        RECT 4.000 88.500 60.550 88.975 ;
        RECT 4.000 88.450 34.675 88.500 ;
      LAYER via ;
        RECT 1.075 91.325 1.350 91.600 ;
        RECT 1.450 91.325 1.725 91.600 ;
        RECT 1.825 91.325 2.100 91.600 ;
        RECT 2.200 91.325 2.475 91.600 ;
        RECT 2.575 91.325 2.850 91.600 ;
        RECT 36.350 90.600 36.700 90.950 ;
        RECT 42.750 90.600 43.100 90.950 ;
        RECT 46.500 90.550 46.900 90.900 ;
        RECT 49.950 90.600 50.300 90.950 ;
        RECT 56.350 90.600 56.700 90.950 ;
        RECT 34.850 89.750 35.200 90.100 ;
        RECT 37.700 89.700 38.050 90.050 ;
        RECT 40.150 90.200 40.500 90.550 ;
        RECT 41.250 89.700 41.600 90.050 ;
        RECT 44.100 89.700 44.450 90.050 ;
        RECT 48.450 89.700 48.850 90.050 ;
        RECT 53.700 90.200 54.050 90.550 ;
        RECT 60.100 90.500 60.450 90.850 ;
        RECT 52.500 89.750 52.850 90.100 ;
        RECT 54.850 89.700 55.200 90.050 ;
        RECT 57.650 89.650 58.000 90.000 ;
        RECT 4.075 88.600 4.350 88.875 ;
        RECT 4.450 88.600 4.725 88.875 ;
        RECT 4.825 88.600 5.100 88.875 ;
        RECT 5.200 88.600 5.475 88.875 ;
        RECT 5.575 88.600 5.850 88.875 ;
      LAYER met2 ;
        RECT 57.600 107.800 58.050 108.300 ;
        RECT 54.750 106.900 55.200 107.400 ;
        RECT 52.500 106.100 52.900 106.500 ;
        RECT 48.400 105.200 48.850 105.700 ;
        RECT 44.050 104.300 44.450 104.800 ;
        RECT 41.300 103.400 41.700 103.900 ;
        RECT 37.700 102.500 38.100 103.000 ;
        RECT 34.850 101.600 35.250 102.100 ;
        RECT 1.000 91.175 3.000 91.750 ;
        RECT 34.900 90.150 35.150 101.600 ;
        RECT 36.300 94.400 36.700 94.900 ;
        RECT 36.350 91.000 36.600 94.400 ;
        RECT 36.300 90.550 36.750 91.000 ;
        RECT 34.800 89.700 35.250 90.150 ;
        RECT 37.750 90.100 38.000 102.500 ;
        RECT 40.100 95.300 40.500 95.800 ;
        RECT 40.150 90.600 40.400 95.300 ;
        RECT 40.100 90.150 40.550 90.600 ;
        RECT 41.350 90.100 41.600 103.400 ;
        RECT 42.750 96.200 43.150 96.700 ;
        RECT 42.800 91.000 43.050 96.200 ;
        RECT 42.700 90.550 43.150 91.000 ;
        RECT 44.150 90.100 44.400 104.300 ;
        RECT 46.500 97.100 46.900 97.600 ;
        RECT 46.550 90.950 46.800 97.100 ;
        RECT 46.450 90.500 46.950 90.950 ;
        RECT 48.500 90.100 48.800 105.200 ;
        RECT 49.950 98.000 50.350 98.500 ;
        RECT 50.000 91.000 50.250 98.000 ;
        RECT 49.900 90.550 50.350 91.000 ;
        RECT 52.600 90.150 52.850 106.100 ;
        RECT 54.850 101.200 55.150 106.900 ;
        RECT 53.700 98.900 54.100 99.400 ;
        RECT 53.750 90.600 54.000 98.900 ;
        RECT 54.860 92.890 55.150 101.200 ;
        RECT 56.350 99.800 56.750 100.300 ;
        RECT 54.850 91.740 55.150 92.890 ;
        RECT 53.650 90.150 54.100 90.600 ;
        RECT 37.650 89.650 38.100 90.100 ;
        RECT 41.200 89.650 41.650 90.100 ;
        RECT 44.050 89.650 44.500 90.100 ;
        RECT 48.400 89.650 48.900 90.100 ;
        RECT 52.450 89.700 52.900 90.150 ;
        RECT 54.890 90.100 55.140 91.740 ;
        RECT 56.400 91.000 56.650 99.800 ;
        RECT 56.300 90.550 56.750 91.000 ;
        RECT 54.800 89.650 55.250 90.100 ;
        RECT 57.700 90.050 57.950 107.800 ;
        RECT 60.100 100.700 60.500 101.200 ;
        RECT 60.150 90.900 60.400 100.700 ;
        RECT 60.050 90.450 60.500 90.900 ;
        RECT 57.600 89.600 58.050 90.050 ;
        RECT 4.000 88.450 6.000 89.025 ;
      LAYER via2 ;
        RECT 57.650 107.850 58.000 108.250 ;
        RECT 54.800 106.950 55.150 107.350 ;
        RECT 52.550 106.150 52.850 106.450 ;
        RECT 48.500 105.250 48.800 105.600 ;
        RECT 44.100 104.400 44.400 104.700 ;
        RECT 41.350 103.450 41.650 103.800 ;
        RECT 37.750 102.600 38.050 102.900 ;
        RECT 34.900 101.700 35.200 102.000 ;
        RECT 1.100 91.325 1.400 91.625 ;
        RECT 1.550 91.325 1.850 91.625 ;
        RECT 2.000 91.325 2.300 91.625 ;
        RECT 2.450 91.325 2.750 91.625 ;
        RECT 36.350 94.500 36.650 94.800 ;
        RECT 40.150 95.400 40.450 95.700 ;
        RECT 42.800 96.300 43.100 96.600 ;
        RECT 46.550 97.200 46.850 97.500 ;
        RECT 50.000 98.100 50.300 98.400 ;
        RECT 53.750 99.000 54.050 99.300 ;
        RECT 56.400 99.900 56.700 100.200 ;
        RECT 60.150 100.800 60.450 101.100 ;
        RECT 4.100 88.600 4.400 88.900 ;
        RECT 4.550 88.600 4.850 88.900 ;
        RECT 5.000 88.600 5.300 88.900 ;
        RECT 5.450 88.600 5.750 88.900 ;
      LAYER met3 ;
        RECT 4.000 108.700 80.500 109.200 ;
        RECT 30.400 107.800 80.500 108.300 ;
        RECT 30.400 106.900 80.500 107.400 ;
        RECT 30.400 106.100 80.500 106.500 ;
        RECT 30.400 105.200 80.500 105.700 ;
        RECT 30.400 104.300 80.500 104.800 ;
        RECT 30.400 103.400 80.500 103.900 ;
        RECT 30.400 102.500 80.500 103.000 ;
        RECT 30.400 101.600 80.500 102.100 ;
        RECT 30.400 100.700 80.500 101.200 ;
        RECT 30.400 99.800 80.500 100.300 ;
        RECT 30.400 98.900 80.500 99.400 ;
        RECT 30.400 98.000 80.500 98.500 ;
        RECT 30.400 97.100 80.500 97.600 ;
        RECT 30.400 96.200 80.500 96.700 ;
        RECT 30.400 95.300 80.500 95.800 ;
        RECT 30.400 94.400 80.500 94.900 ;
        RECT 30.400 93.500 147.000 94.000 ;
        RECT 1.000 91.175 3.000 91.750 ;
        RECT 4.000 88.450 6.000 89.025 ;
      LAYER via3 ;
        RECT 4.050 108.750 4.375 109.125 ;
        RECT 4.475 108.750 4.800 109.125 ;
        RECT 4.900 108.750 5.225 109.125 ;
        RECT 5.325 108.750 5.650 109.125 ;
        RECT 30.650 108.750 31.000 109.150 ;
        RECT 33.400 108.750 33.750 109.150 ;
        RECT 36.150 108.750 36.500 109.150 ;
        RECT 38.900 108.750 39.250 109.150 ;
        RECT 41.700 108.750 42.050 109.150 ;
        RECT 44.450 108.750 44.800 109.150 ;
        RECT 47.200 108.750 47.550 109.150 ;
        RECT 49.950 108.750 50.300 109.150 ;
        RECT 52.700 108.750 53.050 109.150 ;
        RECT 55.500 108.750 55.850 109.150 ;
        RECT 58.250 108.750 58.600 109.150 ;
        RECT 61.000 108.750 61.350 109.150 ;
        RECT 63.750 108.750 64.100 109.150 ;
        RECT 66.500 108.750 66.850 109.150 ;
        RECT 69.300 108.750 69.650 109.150 ;
        RECT 72.050 108.750 72.400 109.150 ;
        RECT 74.800 100.750 75.150 101.150 ;
        RECT 77.550 99.850 77.900 100.250 ;
        RECT 80.300 98.950 80.500 99.350 ;
        RECT 1.075 91.300 1.425 91.650 ;
        RECT 1.525 91.300 1.875 91.650 ;
        RECT 1.975 91.300 2.325 91.650 ;
        RECT 2.425 91.300 2.775 91.650 ;
        RECT 4.075 88.575 4.425 88.925 ;
        RECT 4.525 88.575 4.875 88.925 ;
        RECT 4.975 88.575 5.325 88.925 ;
        RECT 5.425 88.575 5.775 88.925 ;
      LAYER met4 ;
        RECT 30.600 110.520 30.670 110.600 ;
        RECT 30.970 110.520 31.000 110.600 ;
        RECT 30.600 109.200 31.000 110.520 ;
        RECT 33.400 110.520 33.430 110.550 ;
        RECT 33.730 110.520 33.750 110.550 ;
        RECT 33.400 109.200 33.750 110.520 ;
        RECT 36.150 110.520 36.190 110.550 ;
        RECT 36.490 110.520 36.500 110.550 ;
        RECT 36.150 109.200 36.500 110.520 ;
        RECT 38.900 110.520 38.950 110.600 ;
        RECT 41.700 110.520 41.710 110.600 ;
        RECT 42.010 110.520 42.050 110.600 ;
        RECT 38.900 109.200 39.250 110.520 ;
        RECT 41.700 109.200 42.050 110.520 ;
        RECT 44.450 110.520 44.470 110.600 ;
        RECT 44.770 110.520 44.800 110.600 ;
        RECT 44.450 109.200 44.800 110.520 ;
        RECT 47.200 110.520 47.230 110.600 ;
        RECT 47.530 110.520 47.550 110.600 ;
        RECT 47.200 109.200 47.550 110.520 ;
        RECT 49.950 110.520 49.990 110.600 ;
        RECT 50.290 110.520 50.300 110.600 ;
        RECT 49.950 109.200 50.300 110.520 ;
        RECT 52.700 110.520 52.750 110.600 ;
        RECT 55.500 110.520 55.510 110.600 ;
        RECT 55.810 110.520 55.850 110.600 ;
        RECT 52.700 109.200 53.050 110.520 ;
        RECT 55.500 109.200 55.850 110.520 ;
        RECT 58.250 110.520 58.270 110.600 ;
        RECT 58.570 110.520 58.600 110.600 ;
        RECT 58.250 109.200 58.600 110.520 ;
        RECT 61.000 110.520 61.030 110.600 ;
        RECT 61.330 110.520 61.350 110.600 ;
        RECT 61.000 109.200 61.350 110.520 ;
        RECT 63.750 110.520 63.790 110.550 ;
        RECT 64.090 110.520 64.100 110.550 ;
        RECT 63.750 109.200 64.100 110.520 ;
        RECT 66.500 110.520 66.550 110.600 ;
        RECT 69.300 110.520 69.310 110.600 ;
        RECT 69.610 110.520 69.650 110.600 ;
        RECT 66.500 109.200 66.850 110.520 ;
        RECT 69.300 109.200 69.650 110.520 ;
        RECT 72.050 110.520 72.070 110.600 ;
        RECT 72.370 110.520 72.400 110.600 ;
        RECT 72.050 109.200 72.400 110.520 ;
        RECT 74.800 110.520 74.830 110.600 ;
        RECT 75.130 110.520 75.150 110.600 ;
        RECT 30.550 108.700 31.050 109.200 ;
        RECT 33.300 108.700 33.800 109.200 ;
        RECT 36.050 108.700 36.550 109.200 ;
        RECT 38.800 108.700 39.300 109.200 ;
        RECT 41.600 108.700 42.100 109.200 ;
        RECT 44.350 108.700 44.850 109.200 ;
        RECT 47.100 108.700 47.600 109.200 ;
        RECT 49.850 108.700 50.350 109.200 ;
        RECT 52.600 108.700 53.100 109.200 ;
        RECT 55.400 108.700 55.900 109.200 ;
        RECT 58.150 108.700 58.650 109.200 ;
        RECT 60.900 108.700 61.400 109.200 ;
        RECT 63.650 108.700 64.150 109.200 ;
        RECT 66.400 108.700 66.900 109.200 ;
        RECT 69.200 108.700 69.700 109.200 ;
        RECT 71.950 108.700 72.450 109.200 ;
        RECT 74.800 101.200 75.150 110.520 ;
        RECT 77.550 110.520 77.590 110.600 ;
        RECT 77.890 110.520 77.900 110.600 ;
        RECT 74.750 100.700 75.200 101.200 ;
        RECT 77.550 100.300 77.900 110.520 ;
        RECT 80.300 110.520 80.350 110.600 ;
        RECT 77.500 99.800 77.950 100.300 ;
        RECT 80.300 99.400 80.500 110.520 ;
        RECT 80.250 98.900 80.500 99.400 ;
  END
END tt_um_pg_4_bit
END LIBRARY

