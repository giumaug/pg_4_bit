magic
tech sky130A
magscale 1 2
timestamp 1738068025
<< metal1 >>
rect 200 18320 6940 18350
rect 200 18265 215 18320
rect 270 18265 290 18320
rect 345 18265 365 18320
rect 420 18265 440 18320
rect 495 18265 515 18320
rect 570 18265 6940 18320
rect 200 18235 6940 18265
rect 7260 18190 7350 18200
rect 7260 18120 7270 18190
rect 7340 18120 7350 18190
rect 8540 18190 8630 18200
rect 9980 18190 10070 18200
rect 8540 18120 8550 18190
rect 8620 18120 8630 18190
rect 7260 18110 7350 18120
rect 8020 18110 8110 18120
rect 8540 18110 8630 18120
rect 9290 18180 9390 18190
rect 9290 18110 9300 18180
rect 9380 18110 9390 18180
rect 9980 18120 9990 18190
rect 10060 18120 10070 18190
rect 11260 18190 11350 18200
rect 11260 18120 11270 18190
rect 11340 18120 11350 18190
rect 9980 18110 10070 18120
rect 10730 18110 10820 18120
rect 11260 18110 11350 18120
rect 12010 18170 12100 18180
rect 7030 18030 7050 18070
rect 8020 18040 8030 18110
rect 8100 18040 8110 18110
rect 9290 18100 9390 18110
rect 8020 18030 8110 18040
rect 10730 18040 10740 18110
rect 10810 18040 10820 18110
rect 12010 18100 12020 18170
rect 12090 18100 12100 18170
rect 12010 18090 12100 18100
rect 10730 18030 10820 18040
rect 6960 18020 7050 18030
rect 10490 18020 10580 18030
rect 6960 17950 6970 18020
rect 7040 17950 7050 18020
rect 6960 17940 7050 17950
rect 7530 18010 7620 18020
rect 7530 17940 7540 18010
rect 7610 17940 7620 18010
rect 7530 17930 7620 17940
rect 8240 18010 8330 18020
rect 8240 17940 8250 18010
rect 8320 17940 8330 18010
rect 8240 17930 8330 17940
rect 8810 18010 8900 18020
rect 8810 17940 8820 18010
rect 8890 17940 8900 18010
rect 8810 17930 8900 17940
rect 9680 18010 9770 18020
rect 9680 17940 9690 18010
rect 9680 17930 9770 17940
rect 10490 17950 10500 18020
rect 10570 17950 10580 18020
rect 10490 17940 10580 17950
rect 10960 18010 11050 18020
rect 10960 17940 10970 18010
rect 11040 17940 11050 18010
rect 8810 17900 8830 17930
rect 8890 17890 8900 17930
rect 10490 17900 10510 17940
rect 10960 17930 11050 17940
rect 11520 18000 11610 18020
rect 11520 17930 11530 18000
rect 11600 17930 11610 18000
rect 11520 17900 11550 17930
rect 11590 17890 11610 17930
rect 800 17775 6935 17805
rect 800 17720 815 17775
rect 870 17720 890 17775
rect 945 17720 965 17775
rect 1020 17720 1040 17775
rect 1095 17720 1115 17775
rect 1170 17720 6935 17775
rect 800 17690 6935 17720
<< via1 >>
rect 215 18265 270 18320
rect 290 18265 345 18320
rect 365 18265 420 18320
rect 440 18265 495 18320
rect 515 18265 570 18320
rect 7270 18120 7340 18190
rect 8550 18120 8620 18190
rect 9300 18110 9380 18180
rect 9990 18120 10060 18190
rect 11270 18120 11340 18190
rect 8030 18040 8100 18110
rect 10740 18040 10810 18110
rect 12020 18100 12090 18170
rect 6970 17950 7040 18020
rect 7540 17940 7610 18010
rect 8250 17940 8320 18010
rect 8820 17940 8890 18010
rect 9690 17940 9770 18010
rect 10500 17950 10570 18020
rect 10970 17940 11040 18010
rect 11530 17930 11600 18000
rect 815 17720 870 17775
rect 890 17720 945 17775
rect 965 17720 1020 17775
rect 1040 17720 1095 17775
rect 1115 17720 1170 17775
<< metal2 >>
rect 11520 21650 11610 21660
rect 11520 21570 11530 21650
rect 11600 21570 11610 21650
rect 11520 21560 11610 21570
rect 10950 21470 11040 21480
rect 10950 21390 10960 21470
rect 11030 21390 11040 21470
rect 10950 21380 11040 21390
rect 10500 21290 10580 21300
rect 10500 21230 10510 21290
rect 10570 21230 10580 21290
rect 10500 21220 10580 21230
rect 9680 21120 9770 21140
rect 9680 21050 9700 21120
rect 9760 21050 9770 21120
rect 9680 21040 9770 21050
rect 8810 20940 8890 20960
rect 8810 20880 8820 20940
rect 8880 20880 8890 20940
rect 8810 20860 8890 20880
rect 8260 20760 8340 20780
rect 8260 20690 8270 20760
rect 8330 20690 8340 20760
rect 8260 20680 8340 20690
rect 7540 20580 7620 20600
rect 7540 20520 7550 20580
rect 7610 20520 7620 20580
rect 7540 20500 7620 20520
rect 6970 20400 7050 20420
rect 6970 20340 6980 20400
rect 7040 20340 7050 20400
rect 6970 20320 7050 20340
rect 200 18325 600 18350
rect 200 18320 220 18325
rect 280 18320 310 18325
rect 370 18320 400 18325
rect 460 18320 490 18325
rect 550 18320 600 18325
rect 200 18265 215 18320
rect 280 18265 290 18320
rect 570 18265 600 18320
rect 200 18235 600 18265
rect 6980 18030 7030 20320
rect 7260 18960 7340 18980
rect 7260 18900 7270 18960
rect 7330 18900 7340 18960
rect 7260 18880 7340 18900
rect 7270 18200 7320 18880
rect 7260 18190 7350 18200
rect 7260 18120 7270 18190
rect 7340 18120 7350 18190
rect 7260 18110 7350 18120
rect 6960 18020 7050 18030
rect 7550 18020 7600 20500
rect 8020 19140 8100 19160
rect 8020 19080 8030 19140
rect 8090 19080 8100 19140
rect 8020 19060 8100 19080
rect 8030 18120 8080 19060
rect 8020 18110 8110 18120
rect 8020 18040 8030 18110
rect 8100 18040 8110 18110
rect 8020 18030 8110 18040
rect 8270 18020 8320 20680
rect 8550 19320 8630 19340
rect 8550 19260 8560 19320
rect 8620 19260 8630 19320
rect 8550 19240 8630 19260
rect 8560 18200 8610 19240
rect 8540 18190 8630 18200
rect 8540 18120 8550 18190
rect 8620 18120 8630 18190
rect 8540 18110 8630 18120
rect 8830 18020 8880 20860
rect 9300 19500 9380 19520
rect 9300 19440 9310 19500
rect 9370 19440 9380 19500
rect 9300 19420 9380 19440
rect 9310 18190 9360 19420
rect 9290 18180 9390 18190
rect 9290 18110 9300 18180
rect 9380 18110 9390 18180
rect 9290 18100 9390 18110
rect 9700 18020 9760 21040
rect 9990 19680 10070 19700
rect 9990 19620 10000 19680
rect 10060 19620 10070 19680
rect 9990 19600 10070 19620
rect 10000 18200 10050 19600
rect 9980 18190 10070 18200
rect 9980 18120 9990 18190
rect 10060 18120 10070 18190
rect 9980 18110 10070 18120
rect 10520 18030 10570 21220
rect 10970 20240 11030 21380
rect 10740 19860 10820 19880
rect 10740 19800 10750 19860
rect 10810 19800 10820 19860
rect 10740 19780 10820 19800
rect 10750 18120 10800 19780
rect 10972 18578 11030 20240
rect 11270 20040 11350 20060
rect 11270 19980 11280 20040
rect 11340 19980 11350 20040
rect 11270 19960 11350 19980
rect 10970 18348 11030 18578
rect 10730 18110 10820 18120
rect 10730 18040 10740 18110
rect 10810 18040 10820 18110
rect 10730 18030 10820 18040
rect 10490 18020 10580 18030
rect 10978 18020 11028 18348
rect 11280 18200 11330 19960
rect 11260 18190 11350 18200
rect 11260 18120 11270 18190
rect 11340 18120 11350 18190
rect 11260 18110 11350 18120
rect 6960 17950 6970 18020
rect 7040 17950 7050 18020
rect 6960 17940 7050 17950
rect 7530 18010 7620 18020
rect 7530 17940 7540 18010
rect 7610 17940 7620 18010
rect 7530 17930 7620 17940
rect 8240 18010 8330 18020
rect 8240 17940 8250 18010
rect 8320 17940 8330 18010
rect 8240 17930 8330 17940
rect 8810 18010 8900 18020
rect 8810 17940 8820 18010
rect 8890 17940 8900 18010
rect 8810 17930 8900 17940
rect 9680 18010 9780 18020
rect 9680 17940 9690 18010
rect 9770 17940 9780 18010
rect 10490 17950 10500 18020
rect 10570 17950 10580 18020
rect 10490 17940 10580 17950
rect 10960 18010 11050 18020
rect 11540 18010 11590 21560
rect 12020 20220 12100 20240
rect 12020 20160 12030 20220
rect 12090 20160 12100 20220
rect 12020 20140 12100 20160
rect 12030 18180 12080 20140
rect 12010 18170 12100 18180
rect 12010 18100 12020 18170
rect 12090 18100 12100 18170
rect 12010 18090 12100 18100
rect 10960 17940 10970 18010
rect 11040 17940 11050 18010
rect 9680 17930 9780 17940
rect 10960 17930 11050 17940
rect 11520 18000 11610 18010
rect 11520 17930 11530 18000
rect 11600 17930 11610 18000
rect 11520 17920 11610 17930
rect 800 17780 1200 17805
rect 800 17775 820 17780
rect 880 17775 910 17780
rect 970 17775 1000 17780
rect 1060 17775 1090 17780
rect 1150 17775 1200 17780
rect 800 17720 815 17775
rect 880 17720 890 17775
rect 1170 17720 1200 17775
rect 800 17690 1200 17720
<< via2 >>
rect 11530 21570 11600 21650
rect 10960 21390 11030 21470
rect 10510 21230 10570 21290
rect 9700 21050 9760 21120
rect 8820 20880 8880 20940
rect 8270 20690 8330 20760
rect 7550 20520 7610 20580
rect 6980 20340 7040 20400
rect 220 18320 280 18325
rect 310 18320 370 18325
rect 400 18320 460 18325
rect 490 18320 550 18325
rect 220 18265 270 18320
rect 270 18265 280 18320
rect 310 18265 345 18320
rect 345 18265 365 18320
rect 365 18265 370 18320
rect 400 18265 420 18320
rect 420 18265 440 18320
rect 440 18265 460 18320
rect 490 18265 495 18320
rect 495 18265 515 18320
rect 515 18265 550 18320
rect 7270 18900 7330 18960
rect 8030 19080 8090 19140
rect 8560 19260 8620 19320
rect 9310 19440 9370 19500
rect 10000 19620 10060 19680
rect 10750 19800 10810 19860
rect 11280 19980 11340 20040
rect 12030 20160 12090 20220
rect 820 17775 880 17780
rect 910 17775 970 17780
rect 1000 17775 1060 17780
rect 1090 17775 1150 17780
rect 820 17720 870 17775
rect 870 17720 880 17775
rect 910 17720 945 17775
rect 945 17720 965 17775
rect 965 17720 970 17775
rect 1000 17720 1020 17775
rect 1020 17720 1040 17775
rect 1040 17720 1060 17775
rect 1090 17720 1095 17775
rect 1095 17720 1115 17775
rect 1115 17720 1150 17775
<< metal3 >>
rect 800 21830 29400 21840
rect 800 21825 6130 21830
rect 800 21750 810 21825
rect 875 21750 895 21825
rect 960 21750 980 21825
rect 1045 21750 1065 21825
rect 1130 21750 6130 21825
rect 6200 21750 6680 21830
rect 6750 21750 7230 21830
rect 7300 21750 7780 21830
rect 7850 21750 8340 21830
rect 8410 21750 8890 21830
rect 8960 21750 9440 21830
rect 9510 21750 9990 21830
rect 10060 21750 10540 21830
rect 10610 21750 11100 21830
rect 11170 21750 11650 21830
rect 11720 21750 12200 21830
rect 12270 21750 12750 21830
rect 12820 21750 13300 21830
rect 13370 21750 13860 21830
rect 13930 21750 14410 21830
rect 14480 21750 29400 21830
rect 800 21740 29400 21750
rect 6080 21650 29400 21660
rect 6080 21570 11530 21650
rect 11600 21570 23780 21650
rect 23860 21570 29400 21650
rect 6080 21560 29400 21570
rect 6080 21470 29400 21480
rect 6080 21390 10960 21470
rect 11030 21390 24340 21470
rect 24410 21390 29400 21470
rect 6080 21380 29400 21390
rect 24880 21300 24990 21310
rect 6080 21290 24880 21300
rect 6080 21230 10510 21290
rect 10570 21230 24880 21290
rect 6080 21220 24880 21230
rect 24980 21220 29400 21300
rect 24880 21210 24990 21220
rect 6080 21130 29400 21140
rect 6080 21120 25450 21130
rect 6080 21050 9700 21120
rect 9760 21050 25450 21120
rect 6080 21048 25450 21050
rect 25530 21048 29400 21130
rect 6080 21040 29400 21048
rect 6080 20950 29400 20960
rect 6080 20940 26000 20950
rect 6080 20880 8820 20940
rect 8880 20880 26000 20940
rect 6080 20870 26000 20880
rect 26080 20870 29400 20950
rect 6080 20860 29400 20870
rect 6080 20770 29400 20780
rect 6080 20760 26540 20770
rect 6080 20690 8270 20760
rect 8330 20690 26540 20760
rect 26620 20690 29400 20770
rect 6080 20680 29400 20690
rect 6080 20590 29400 20600
rect 6080 20580 27100 20590
rect 6080 20520 7550 20580
rect 7610 20520 27100 20580
rect 6080 20510 27100 20520
rect 27180 20510 29400 20590
rect 6080 20500 29400 20510
rect 6080 20410 29400 20420
rect 6080 20400 27640 20410
rect 6080 20340 6980 20400
rect 7040 20340 27640 20400
rect 6080 20330 27640 20340
rect 27720 20330 29400 20410
rect 6080 20320 29400 20330
rect 6080 20230 29400 20240
rect 6080 20220 14960 20230
rect 6080 20160 12030 20220
rect 12090 20160 14960 20220
rect 6080 20150 14960 20160
rect 15030 20150 29400 20230
rect 6080 20140 29400 20150
rect 6080 20050 29400 20060
rect 6080 20040 15510 20050
rect 6080 19980 11280 20040
rect 11340 19980 15510 20040
rect 6080 19970 15510 19980
rect 15580 19970 29400 20050
rect 6080 19960 29400 19970
rect 6080 19870 29400 19880
rect 6080 19860 16060 19870
rect 6080 19800 10750 19860
rect 10810 19800 16060 19860
rect 6080 19790 16060 19800
rect 16130 19790 29400 19870
rect 6080 19780 29400 19790
rect 6080 19690 29400 19700
rect 6080 19680 16620 19690
rect 6080 19620 10000 19680
rect 10060 19620 16620 19680
rect 6080 19610 16620 19620
rect 16690 19610 29400 19690
rect 6080 19600 29400 19610
rect 6080 19510 29400 19520
rect 6080 19500 17160 19510
rect 6080 19440 9310 19500
rect 9370 19440 17160 19500
rect 6080 19430 17160 19440
rect 17240 19430 29400 19510
rect 6080 19420 29400 19430
rect 6080 19330 29400 19340
rect 6080 19320 17720 19330
rect 6080 19260 8560 19320
rect 8620 19260 17720 19320
rect 6080 19250 17720 19260
rect 17800 19250 29400 19330
rect 6080 19240 29400 19250
rect 6080 19150 29400 19160
rect 6080 19140 18260 19150
rect 6080 19080 8030 19140
rect 8090 19080 18260 19140
rect 6080 19070 18260 19080
rect 18340 19070 29400 19150
rect 6080 19060 29400 19070
rect 6080 18970 29400 18980
rect 6080 18960 18820 18970
rect 6080 18900 7270 18960
rect 7330 18900 18820 18960
rect 6080 18890 18820 18900
rect 18900 18890 29400 18970
rect 6080 18880 29400 18890
rect 6080 18700 29400 18800
rect 200 18330 600 18350
rect 200 18260 215 18330
rect 285 18260 305 18330
rect 375 18260 395 18330
rect 465 18260 485 18330
rect 555 18260 600 18330
rect 200 18235 600 18260
rect 800 17785 1200 17805
rect 800 17715 815 17785
rect 885 17715 905 17785
rect 975 17715 995 17785
rect 1065 17715 1085 17785
rect 1155 17715 1200 17785
rect 800 17690 1200 17715
<< via3 >>
rect 810 21750 875 21825
rect 895 21750 960 21825
rect 980 21750 1045 21825
rect 1065 21750 1130 21825
rect 6130 21750 6200 21830
rect 6680 21750 6750 21830
rect 7230 21750 7300 21830
rect 7780 21750 7850 21830
rect 8340 21750 8410 21830
rect 8890 21750 8960 21830
rect 9440 21750 9510 21830
rect 9990 21750 10060 21830
rect 10540 21750 10610 21830
rect 11100 21750 11170 21830
rect 11650 21750 11720 21830
rect 12200 21750 12270 21830
rect 12750 21750 12820 21830
rect 13300 21750 13370 21830
rect 13860 21750 13930 21830
rect 14410 21750 14480 21830
rect 23780 21570 23860 21650
rect 24340 21390 24410 21470
rect 24880 21220 24980 21300
rect 25450 21048 25530 21130
rect 26000 20870 26080 20950
rect 26540 20690 26620 20770
rect 27100 20510 27180 20590
rect 27640 20330 27720 20410
rect 14960 20150 15030 20230
rect 15510 19970 15580 20050
rect 16060 19790 16130 19870
rect 16620 19610 16690 19690
rect 17160 19430 17240 19510
rect 17720 19250 17800 19330
rect 18260 19070 18340 19150
rect 18820 18890 18900 18970
rect 215 18325 285 18330
rect 215 18265 220 18325
rect 220 18265 280 18325
rect 280 18265 285 18325
rect 215 18260 285 18265
rect 305 18325 375 18330
rect 305 18265 310 18325
rect 310 18265 370 18325
rect 370 18265 375 18325
rect 305 18260 375 18265
rect 395 18325 465 18330
rect 395 18265 400 18325
rect 400 18265 460 18325
rect 460 18265 465 18325
rect 395 18260 465 18265
rect 485 18325 555 18330
rect 485 18265 490 18325
rect 490 18265 550 18325
rect 550 18265 555 18325
rect 485 18260 555 18265
rect 815 17780 885 17785
rect 815 17720 820 17780
rect 820 17720 880 17780
rect 880 17720 885 17780
rect 815 17715 885 17720
rect 905 17780 975 17785
rect 905 17720 910 17780
rect 910 17720 970 17780
rect 970 17720 975 17780
rect 905 17715 975 17720
rect 995 17780 1065 17785
rect 995 17720 1000 17780
rect 1000 17720 1060 17780
rect 1060 17720 1065 17780
rect 995 17715 1065 17720
rect 1085 17780 1155 17785
rect 1085 17720 1090 17780
rect 1090 17720 1150 17780
rect 1150 17720 1155 17780
rect 1085 17715 1155 17720
<< metal4 >>
rect 200 18330 600 44152
rect 200 18260 215 18330
rect 285 18260 305 18330
rect 375 18260 395 18330
rect 465 18260 485 18330
rect 555 18260 600 18330
rect 200 1000 600 18260
rect 800 21825 1200 44152
rect 6134 22120 6194 22304
rect 6120 21840 6200 22120
rect 6686 22110 6746 22304
rect 7238 22110 7298 22304
rect 7790 22120 7850 22304
rect 8342 22120 8402 22304
rect 8894 22120 8954 22304
rect 9446 22120 9506 22304
rect 9998 22120 10058 22304
rect 10550 22120 10610 22304
rect 11102 22120 11162 22304
rect 11654 22120 11714 22304
rect 12206 22120 12266 22304
rect 6680 21840 6750 22110
rect 7230 21840 7300 22110
rect 7780 21840 7850 22120
rect 8340 21840 8410 22120
rect 8890 21840 8960 22120
rect 9440 21840 9510 22120
rect 9990 21840 10060 22120
rect 10540 21840 10610 22120
rect 11100 21840 11170 22120
rect 11650 21840 11720 22120
rect 12200 21840 12270 22120
rect 12758 22110 12818 22304
rect 13310 22120 13370 22304
rect 13862 22120 13922 22304
rect 14414 22120 14474 22304
rect 14966 22120 15026 22304
rect 15518 22120 15578 22304
rect 16070 22120 16130 22304
rect 16622 22120 16682 22304
rect 17174 22120 17234 22304
rect 17726 22120 17786 22304
rect 18278 22120 18338 22304
rect 18830 22120 18890 22304
rect 12750 21840 12820 22110
rect 13300 21840 13370 22120
rect 13860 21840 13930 22120
rect 14410 21840 14480 22120
rect 800 21750 810 21825
rect 875 21750 895 21825
rect 960 21750 980 21825
rect 1045 21750 1065 21825
rect 1130 21750 1200 21825
rect 800 17785 1200 21750
rect 6110 21830 6210 21840
rect 6110 21750 6130 21830
rect 6200 21750 6210 21830
rect 6110 21740 6210 21750
rect 6660 21830 6760 21840
rect 6660 21750 6680 21830
rect 6750 21750 6760 21830
rect 6660 21740 6760 21750
rect 7210 21830 7310 21840
rect 7210 21750 7230 21830
rect 7300 21750 7310 21830
rect 7210 21740 7310 21750
rect 7760 21830 7860 21840
rect 7760 21750 7780 21830
rect 7850 21750 7860 21830
rect 7760 21740 7860 21750
rect 8320 21830 8420 21840
rect 8320 21750 8340 21830
rect 8410 21750 8420 21830
rect 8320 21740 8420 21750
rect 8870 21830 8970 21840
rect 8870 21750 8890 21830
rect 8960 21750 8970 21830
rect 8870 21740 8970 21750
rect 9420 21830 9520 21840
rect 9420 21750 9440 21830
rect 9510 21750 9520 21830
rect 9420 21740 9520 21750
rect 9970 21830 10070 21840
rect 9970 21750 9990 21830
rect 10060 21750 10070 21830
rect 9970 21740 10070 21750
rect 10520 21830 10620 21840
rect 10520 21750 10540 21830
rect 10610 21750 10620 21830
rect 10520 21740 10620 21750
rect 11080 21830 11180 21840
rect 11080 21750 11100 21830
rect 11170 21750 11180 21830
rect 11080 21740 11180 21750
rect 11630 21830 11730 21840
rect 11630 21750 11650 21830
rect 11720 21750 11730 21830
rect 11630 21740 11730 21750
rect 12180 21830 12280 21840
rect 12180 21750 12200 21830
rect 12270 21750 12280 21830
rect 12180 21740 12280 21750
rect 12730 21830 12830 21840
rect 12730 21750 12750 21830
rect 12820 21750 12830 21830
rect 12730 21740 12830 21750
rect 13280 21830 13380 21840
rect 13280 21750 13300 21830
rect 13370 21750 13380 21830
rect 13280 21740 13380 21750
rect 13840 21830 13940 21840
rect 13840 21750 13860 21830
rect 13930 21750 13940 21830
rect 13840 21740 13940 21750
rect 14390 21830 14490 21840
rect 14390 21750 14410 21830
rect 14480 21750 14490 21830
rect 14390 21740 14490 21750
rect 14960 20240 15030 22120
rect 14950 20230 15040 20240
rect 14950 20150 14960 20230
rect 15030 20150 15040 20230
rect 14950 20140 15040 20150
rect 15510 20060 15580 22120
rect 15500 20050 15590 20060
rect 15500 19970 15510 20050
rect 15580 19970 15590 20050
rect 15500 19960 15590 19970
rect 16060 19880 16130 22120
rect 16050 19870 16140 19880
rect 16050 19790 16060 19870
rect 16130 19790 16140 19870
rect 16050 19780 16140 19790
rect 16620 19700 16690 22120
rect 16610 19690 16700 19700
rect 16610 19610 16620 19690
rect 16690 19610 16700 19690
rect 16610 19600 16700 19610
rect 17160 19520 17240 22120
rect 17150 19510 17250 19520
rect 17150 19430 17160 19510
rect 17240 19430 17250 19510
rect 17150 19420 17250 19430
rect 17720 19340 17800 22120
rect 17710 19330 17810 19340
rect 17710 19250 17720 19330
rect 17800 19250 17810 19330
rect 17710 19240 17810 19250
rect 18260 19160 18340 22120
rect 18250 19150 18350 19160
rect 18250 19070 18260 19150
rect 18340 19070 18350 19150
rect 18250 19060 18350 19070
rect 18820 18980 18900 22120
rect 19382 22104 19442 22304
rect 19934 22104 19994 22304
rect 20486 22104 20546 22304
rect 21038 22104 21098 22304
rect 21590 22104 21650 22304
rect 22142 22104 22202 22304
rect 22694 22104 22754 22304
rect 23246 22104 23306 22304
rect 23798 22120 23858 22304
rect 23790 21660 23860 22120
rect 23770 21650 23870 21660
rect 23770 21570 23780 21650
rect 23860 21570 23870 21650
rect 23770 21560 23870 21570
rect 24350 21480 24410 22304
rect 24902 22120 24962 22304
rect 25454 22130 25514 22304
rect 24330 21470 24420 21480
rect 24330 21390 24340 21470
rect 24410 21390 24420 21470
rect 24330 21380 24420 21390
rect 24900 21310 24970 22120
rect 24870 21300 24990 21310
rect 24870 21220 24880 21300
rect 24980 21220 24990 21300
rect 24870 21210 24990 21220
rect 25450 21140 25530 22130
rect 26006 22120 26066 22304
rect 26558 22120 26618 22304
rect 27110 22120 27170 22304
rect 27662 22170 27722 22304
rect 25430 21130 25540 21140
rect 25430 21048 25450 21130
rect 25530 21048 25540 21130
rect 25430 21040 25540 21048
rect 26000 20960 26080 22120
rect 25980 20950 26090 20960
rect 25980 20870 26000 20950
rect 26080 20870 26090 20950
rect 25980 20860 26090 20870
rect 26540 20780 26620 22120
rect 26520 20770 26630 20780
rect 26520 20690 26540 20770
rect 26620 20690 26630 20770
rect 26520 20680 26630 20690
rect 27100 20600 27180 22120
rect 27640 22104 27722 22170
rect 28214 22104 28274 22304
rect 28766 22104 28826 22304
rect 29318 22104 29378 22304
rect 27080 20590 27190 20600
rect 27080 20510 27100 20590
rect 27180 20510 27190 20590
rect 27080 20500 27190 20510
rect 27640 20420 27720 22104
rect 27620 20410 27730 20420
rect 27620 20330 27640 20410
rect 27720 20330 27730 20410
rect 27620 20320 27730 20330
rect 18810 18970 18910 18980
rect 18810 18890 18820 18970
rect 18900 18890 18910 18970
rect 18810 18880 18910 18890
rect 800 17715 815 17785
rect 885 17715 905 17785
rect 975 17715 995 17785
rect 1065 17715 1085 17785
rect 1155 17715 1200 17785
rect 800 1000 1200 17715
use adder_1  adder_1_0
timestamp 1700079872
transform 1 0 6960 0 1 17750
box -80 -50 5188 590
<< labels >>
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 200 1000 600 44152 1 FreeSans 4 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 4 0 0 0 VGND
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32972800 22839296
<< end >>
