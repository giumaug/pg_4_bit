magic
tech sky130A
magscale 1 2
timestamp 1700079872
<< nwell >>
rect 433 259 473 580
rect 1184 259 1204 580
rect 1207 259 1247 579
rect 1724 259 1754 580
rect 3167 259 3191 580
rect 3900 259 3921 580
rect 4446 259 4474 580
<< pwell >>
rect 343 45 523 200
rect 1148 45 1278 183
rect 1619 46 1802 200
rect 2422 45 2522 193
rect 2590 46 2713 183
rect 3061 45 3244 200
rect 3863 46 3994 183
rect 4369 46 4519 201
<< locali >>
rect 412 525 444 559
rect 480 525 513 559
rect 1144 525 1180 559
rect 1215 525 1245 559
rect 1693 525 1724 559
rect 1760 525 1793 559
rect 2428 525 2450 559
rect 2485 525 2512 559
rect 2592 525 2625 559
rect 2660 525 2678 559
rect 3132 525 3163 559
rect 3198 525 3231 559
rect 3862 525 3898 559
rect 3933 525 3962 559
rect 4411 525 4443 559
rect 4478 525 4512 559
rect 340 420 375 454
rect 397 -20 444 15
rect 480 -20 515 15
rect 1147 -19 1174 15
rect 1210 -19 1246 15
rect 1686 -19 1725 15
rect 1760 -19 1795 15
rect 2429 -19 2450 15
rect 2485 -19 2516 15
rect 2592 -19 2620 15
rect 2655 -19 2679 15
rect 3124 -19 3163 15
rect 3198 -19 3229 15
rect 3864 -19 3898 15
rect 3933 -19 3960 15
rect 4405 -19 4443 15
rect 4478 -19 4513 15
<< viali >>
rect 79 525 113 559
rect 444 525 480 559
rect 1180 525 1215 559
rect 1724 525 1760 559
rect 2450 525 2485 559
rect 2625 525 2660 559
rect 3163 525 3198 559
rect 3898 525 3933 559
rect 4443 525 4478 559
rect 325 381 359 415
rect 1605 381 1639 415
rect 2355 373 2389 407
rect 3043 381 3077 415
rect 4323 381 4357 415
rect 5073 373 5107 407
rect 1075 305 1109 339
rect 3793 305 3827 339
rect 32 213 66 247
rect 173 213 207 247
rect 593 213 627 247
rect 710 213 744 247
rect 1312 213 1346 247
rect 1453 213 1487 247
rect 1873 213 1907 247
rect 1990 213 2024 247
rect 2750 213 2784 247
rect 2891 213 2925 247
rect 3428 213 3462 247
rect 3563 213 3597 247
rect 4030 213 4064 247
rect 4171 213 4205 247
rect 4591 213 4625 247
rect 4708 213 4742 247
rect 444 -20 480 15
rect 1174 -19 1210 15
rect 1725 -19 1760 15
rect 2450 -19 2485 15
rect 2620 -19 2655 15
rect 3163 -19 3198 15
rect 3898 -19 3933 15
rect 4443 -19 4478 15
<< metal1 >>
rect 413 559 511 590
rect 413 525 444 559
rect 480 525 511 559
rect 413 494 511 525
rect 1145 559 1242 590
rect 1145 525 1180 559
rect 1215 525 1242 559
rect 1145 494 1242 525
rect 1693 559 1791 590
rect 1693 525 1724 559
rect 1760 525 1791 559
rect 1693 494 1791 525
rect 2425 559 2513 590
rect 2425 525 2450 559
rect 2485 525 2513 559
rect 2425 494 2513 525
rect 2595 559 2684 590
rect 2595 525 2625 559
rect 2660 525 2684 559
rect 2595 494 2684 525
rect 3130 559 3231 590
rect 3130 525 3163 559
rect 3198 525 3231 559
rect 3130 494 3231 525
rect 3864 559 3962 590
rect 3864 525 3898 559
rect 3933 525 3962 559
rect 3864 494 3962 525
rect 4411 559 4512 590
rect 4411 525 4443 559
rect 4478 525 4512 559
rect 4411 494 4512 525
rect 310 415 400 425
rect 310 381 325 415
rect 359 381 400 415
rect 310 375 400 381
rect 1590 415 1680 425
rect 1590 381 1605 415
rect 1639 381 1680 415
rect 1590 375 1680 381
rect 2340 407 2410 425
rect 2340 373 2355 407
rect 2389 373 2410 407
rect 1066 339 1130 370
rect 2340 360 2410 373
rect 3023 415 3113 425
rect 3023 381 3043 415
rect 3077 381 3113 415
rect 3023 369 3113 381
rect 4308 415 4398 425
rect 4308 381 4323 415
rect 4357 381 4398 415
rect 4308 370 4398 381
rect 5058 407 5128 425
rect 5058 373 5073 407
rect 5107 373 5128 407
rect 5058 360 5128 373
rect 20 301 760 330
rect 20 300 634 301
rect 20 247 80 300
rect 20 213 32 247
rect 66 213 80 247
rect 20 200 80 213
rect 160 247 220 260
rect 160 213 173 247
rect 207 213 220 247
rect 160 210 220 213
rect 157 190 220 210
rect 579 247 640 260
rect 579 213 593 247
rect 627 213 640 247
rect 579 190 640 213
rect 690 247 760 301
rect 1066 305 1075 339
rect 1109 305 1130 339
rect 3778 339 3848 355
rect 1066 286 1130 305
rect 1300 300 2040 330
rect 690 213 710 247
rect 744 213 760 247
rect 690 200 760 213
rect 1300 247 1360 300
rect 1300 213 1312 247
rect 1346 213 1360 247
rect 1300 200 1360 213
rect 1440 247 1500 260
rect 1440 213 1453 247
rect 1487 213 1500 247
rect 1440 200 1500 213
rect 1860 247 1930 260
rect 1860 213 1873 247
rect 1907 213 1930 247
rect 157 160 640 190
rect 1440 170 1470 200
rect 1860 170 1930 213
rect 1980 247 2040 300
rect 1980 213 1990 247
rect 2024 213 2040 247
rect 1980 200 2040 213
rect 2738 300 3468 330
rect 2738 247 2798 300
rect 2738 213 2750 247
rect 2784 213 2798 247
rect 2738 200 2798 213
rect 2878 247 2938 260
rect 2878 213 2891 247
rect 2925 213 2938 247
rect 1440 141 1930 170
rect 1500 140 1930 141
rect 2878 170 2938 213
rect 3418 247 3468 300
rect 3778 305 3793 339
rect 3827 305 3848 339
rect 3778 290 3848 305
rect 4018 300 4758 330
rect 3418 213 3428 247
rect 3462 213 3468 247
rect 3418 200 3468 213
rect 3548 247 3608 260
rect 3548 213 3563 247
rect 3597 213 3608 247
rect 3548 170 3608 213
rect 4018 247 4078 300
rect 4018 213 4030 247
rect 4064 213 4078 247
rect 4018 199 4078 213
rect 4158 247 4218 260
rect 4588 259 4638 260
rect 4158 213 4171 247
rect 4205 213 4218 247
rect 2878 140 3608 170
rect 4158 170 4218 213
rect 4578 247 4638 259
rect 4578 213 4591 247
rect 4625 213 4638 247
rect 4578 170 4638 213
rect 4698 247 4758 300
rect 4698 213 4708 247
rect 4742 213 4758 247
rect 4698 200 4758 213
rect 4158 140 4638 170
rect 405 15 515 45
rect 405 -20 444 15
rect 480 -20 515 15
rect 405 -50 515 -20
rect 1144 15 1246 46
rect 1690 15 1796 46
rect 1144 -19 1174 15
rect 1210 -19 1246 15
rect 1686 -19 1725 15
rect 1760 -19 1796 15
rect 1144 -50 1246 -19
rect 1690 -50 1796 -19
rect 2423 15 2513 46
rect 2423 -19 2450 15
rect 2485 -19 2513 15
rect 2423 -50 2513 -19
rect 2599 15 2684 46
rect 2599 -19 2620 15
rect 2655 -19 2684 15
rect 2599 -50 2684 -19
rect 3131 15 3231 46
rect 3131 -19 3163 15
rect 3198 -19 3231 15
rect 3131 -50 3231 -19
rect 3864 15 3962 46
rect 3864 -19 3898 15
rect 3933 -19 3962 15
rect 3864 -50 3962 -19
rect 4410 15 4513 46
rect 4410 -19 4443 15
rect 4478 -19 4513 15
rect 4410 -50 4513 -19
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1691611044
transform 1 0 -42 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1691611044
transform 1 0 1238 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1691611044
transform 1 0 2676 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1691611044
transform 1 0 3956 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 2508 0 1 -2
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 508 0 1 -2
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 1788 0 1 -2
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 3226 0 1 -2
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4506 0 1 -2
box -38 -48 682 592
<< labels >>
flabel metal1 1300 240 1300 240 1 FreeSans 320 0 0 0 A2
port 3 n
flabel viali 610 240 610 240 1 FreeSans 192 0 0 0 B1
port 2 n
flabel viali 1890 242 1890 242 1 FreeSans 192 0 0 0 B2
port 4 n
flabel viali 1090 330 1090 330 1 FreeSans 192 0 0 0 P1
port 10 n
flabel viali 340 405 340 405 1 FreeSans 128 0 0 0 G1
port 9 n
flabel viali 1620 405 1620 405 1 FreeSans 160 0 0 0 G2
port 11 n
flabel viali 2370 400 2370 400 1 FreeSans 128 0 0 0 P2
port 12 n
flabel viali 2768 240 2768 240 1 FreeSans 256 0 0 0 A3
port 5 n
flabel viali 3578 240 3578 240 1 FreeSans 192 0 0 0 B3
port 6 n
flabel viali 4046 240 4046 240 1 FreeSans 192 0 0 0 A4
port 7 n
flabel viali 4610 238 4610 238 1 FreeSans 192 0 0 0 B4
port 8 n
flabel viali 5088 400 5088 400 1 FreeSans 128 0 0 0 P4
port 16 n
flabel viali 3808 326 3808 326 1 FreeSans 256 0 0 0 P3
port 14 n
flabel viali 3058 400 3058 400 1 FreeSans 160 0 0 0 G3
port 13 n
flabel viali 4336 400 4336 400 1 FreeSans 160 0 0 0 G4
port 15 n
flabel metal1 s -30 570 -30 570 1 FreeSans 128 0 0 0 VDD
port 17 n
flabel metal1 s -35 25 -35 25 1 FreeSans 96 0 0 0 GND
port 18 n
flabel space 2548 447 2548 447 1 FreeSans 128 0 0 0 VPB
port 19 n
flabel space 2550 135 2550 135 1 FreeSans 128 0 0 0 VNB
port 20 n
flabel viali 45 230 45 230 1 FreeSans 160 0 0 0 A1
port 1 n
<< end >>
