* NGSPICE file created from adder.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.229 ps=1.57 w=0.65 l=0.15
**devattr s=10270,288 d=3575,185
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5500,255
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=10270,288
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
**devattr s=3575,185 d=3640,186
C0 VGND a_299_297# 0.00772f
C1 B1 X 3.04e-20
C2 VPWR VGND 0.0579f
C3 A2 VPB 0.0373f
C4 VPB A1 0.0264f
C5 A2 a_81_21# 7.47e-19
C6 B1 a_299_297# 0.00863f
C7 a_81_21# A1 0.0568f
C8 a_81_21# a_384_47# 0.00138f
C9 VPWR B1 0.0196f
C10 A2 a_299_297# 0.0468f
C11 a_81_21# VPB 0.0593f
C12 a_299_297# A1 0.0585f
C13 VPWR A2 0.0201f
C14 a_384_47# a_299_297# 1.48e-19
C15 VPWR A1 0.0209f
C16 B1 VGND 0.0181f
C17 X VPB 0.0108f
C18 VPWR a_384_47# 4.08e-19
C19 X a_81_21# 0.112f
C20 a_299_297# VPB 0.0111f
C21 A2 VGND 0.0495f
C22 VPWR VPB 0.068f
C23 a_81_21# a_299_297# 0.0821f
C24 VGND A1 0.0786f
C25 VGND a_384_47# 0.00366f
C26 VPWR a_81_21# 0.146f
C27 VPWR X 0.0847f
C28 B1 A1 0.0817f
C29 VGND VPB 0.00713f
C30 VPWR a_299_297# 0.202f
C31 VGND a_81_21# 0.173f
C32 A2 A1 0.0921f
C33 X VGND 0.0512f
C34 B1 VPB 0.0387f
C35 a_384_47# A1 0.00884f
C36 B1 a_81_21# 0.148f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.139 ps=0.987 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.332 ps=2.35 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.139 ps=0.987 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139 pd=0.987 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139 pd=0.987 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.238 ps=1.62 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
C0 VPB VPWR 0.077f
C1 a_109_47# VGND 0.00223f
C2 D a_27_47# 0.107f
C3 a_303_47# a_27_47# 0.00119f
C4 C D 0.18f
C5 VPB A 0.0907f
C6 a_27_47# a_197_47# 0.00167f
C7 a_303_47# C 0.00527f
C8 B a_27_47# 0.13f
C9 VGND D 0.0898f
C10 a_109_47# VPWR 4.66e-19
C11 C a_197_47# 0.00123f
C12 a_303_47# VGND 0.00381f
C13 C B 0.161f
C14 X D 0.00746f
C15 VGND a_197_47# 0.00387f
C16 B VGND 0.0453f
C17 VPWR D 0.0207f
C18 a_303_47# VPWR 4.83e-19
C19 C a_27_47# 0.0516f
C20 VPWR a_197_47# 5.24e-19
C21 B VPWR 0.0231f
C22 VGND a_27_47# 0.132f
C23 C VGND 0.0408f
C24 A B 0.0839f
C25 X a_27_47# 0.0754f
C26 VPB D 0.0782f
C27 VPWR a_27_47# 0.326f
C28 X VGND 0.0903f
C29 C VPWR 0.021f
C30 A a_27_47# 0.153f
C31 VPB B 0.0643f
C32 VPWR VGND 0.0662f
C33 X VPWR 0.0945f
C34 A VGND 0.0151f
C35 a_109_47# B 0.00153f
C36 VPB a_27_47# 0.082f
C37 a_303_47# D 0.00119f
C38 VPB C 0.0609f
C39 A VPWR 0.044f
C40 VPB VGND 0.00852f
C41 a_109_47# a_27_47# 0.00578f
C42 B a_197_47# 0.00623f
C43 VPB X 0.0111f
C44 a_109_47# C 1.72e-20
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt adder_2 CI P1 G1 P2 G2 P3 G3 P4 G4 CO VDD SUB sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_1/X
+ sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__and4_1_0/a_109_47#
+ sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_3/a_299_297#
+ sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ sky130_fd_sc_hd__a21o_1_3/a_384_47#
Xsky130_fd_sc_hd__a21o_1_0 G1 P2 G2 SUB SUB VDD VDD sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__a21o_1_0/X P3 G3 SUB SUB VDD VDD sky130_fd_sc_hd__a21o_1_1/X
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__a21o_1_1/X P4 G4 SUB SUB VDD VDD sky130_fd_sc_hd__a21o_1_2/X
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_3 sky130_fd_sc_hd__and4_1_0/X CI sky130_fd_sc_hd__a21o_1_2/X
+ SUB SUB VDD VDD CO sky130_fd_sc_hd__a21o_1_3/a_384_47# sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ sky130_fd_sc_hd__a21o_1_3/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__and4_1_0 P4 P2 P3 P1 SUB SUB VDD VDD sky130_fd_sc_hd__and4_1_0/X
+ sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__and4_1_0/a_303_47#
+ sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1
C0 sky130_fd_sc_hd__and4_1_0/X VDD 0.0202f
C1 P4 G4 0.02f
C2 sky130_fd_sc_hd__a21o_1_1/X G4 0.0897f
C3 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__a21o_1_0/X 5.18e-21
C4 sky130_fd_sc_hd__a21o_1_0/X VDD 0.0377f
C5 sky130_fd_sc_hd__and4_1_0/a_197_47# P2 2.63e-19
C6 P2 CO 4.84e-19
C7 CI sky130_fd_sc_hd__a21o_1_2/X 0.00156f
C8 sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__and4_1_0/X 1.78e-19
C9 sky130_fd_sc_hd__and4_1_0/X CO 0.13f
C10 VDD sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00151f
C11 sky130_fd_sc_hd__a21o_1_2/a_299_297# P3 0.00159f
C12 VDD sky130_fd_sc_hd__a21o_1_2/a_384_47# -4.08e-19
C13 sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__a21o_1_0/X 5.93e-21
C14 sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD -0.00647f
C15 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0335f
C16 G3 VDD -6.71e-19
C17 sky130_fd_sc_hd__a21o_1_3/a_81_21# VDD -0.0123f
C18 SUB sky130_fd_sc_hd__a21o_1_1/a_384_47# -1.89e-19
C19 CI sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.00978f
C20 P2 P1 0.0215f
C21 sky130_fd_sc_hd__and4_1_0/a_303_47# P3 4.7e-19
C22 P4 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0108f
C23 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__a21o_1_2/X 4.26e-19
C24 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0193f
C25 P2 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0566f
C26 VDD P3 0.0048f
C27 sky130_fd_sc_hd__and4_1_0/X P1 0.00732f
C28 sky130_fd_sc_hd__a21o_1_2/X VDD 1.21f
C29 P2 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0301f
C30 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_384_47# 0.00135f
C31 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.69e-20
C32 P4 VDD 0.0594f
C33 sky130_fd_sc_hd__a21o_1_1/X VDD 0.0255f
C34 P2 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0456f
C35 VDD G2 0.0175f
C36 sky130_fd_sc_hd__a21o_1_0/X P1 1.23e-20
C37 SUB sky130_fd_sc_hd__and4_1_0/a_109_47# -6.28e-20
C38 VDD G1 0.0196f
C39 VDD sky130_fd_sc_hd__a21o_1_3/a_299_297# -5.68e-32
C40 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.2e-19
C41 sky130_fd_sc_hd__a21o_1_3/a_81_21# CO 0.00936f
C42 sky130_fd_sc_hd__and4_1_0/a_27_47# VDD -0.0199f
C43 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00259f
C44 sky130_fd_sc_hd__and4_1_0/a_197_47# P3 0.0016f
C45 CO P3 0.0012f
C46 G4 VDD -0.00221f
C47 sky130_fd_sc_hd__a21o_1_2/X CO 0.0504f
C48 G3 P1 3.23e-21
C49 sky130_fd_sc_hd__a21o_1_3/a_81_21# P1 0.00196f
C50 P1 P3 0.0581f
C51 sky130_fd_sc_hd__a21o_1_2/X P1 0.0247f
C52 P3 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00415f
C53 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_0/a_384_47# 1.32e-20
C54 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0334f
C55 sky130_fd_sc_hd__and4_1_0/a_27_47# CO 0.00246f
C56 sky130_fd_sc_hd__a21o_1_2/a_81_21# P3 0.0706f
C57 P4 P1 4.35e-19
C58 sky130_fd_sc_hd__a21o_1_1/X P1 4.83e-20
C59 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.02f
C60 sky130_fd_sc_hd__a21o_1_0/a_384_47# G1 4.61e-19
C61 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0338f
C62 P4 sky130_fd_sc_hd__a21o_1_1/a_299_297# 1.23e-19
C63 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.46e-21
C64 CI VDD 0.00996f
C65 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 1.65e-19
C66 VDD sky130_fd_sc_hd__a21o_1_3/a_384_47# -1.62e-19
C67 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0421f
C68 P4 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00149f
C69 P1 sky130_fd_sc_hd__a21o_1_3/a_299_297# 2.61e-19
C70 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0315f
C71 sky130_fd_sc_hd__and4_1_0/a_27_47# P1 0.019f
C72 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 6.97e-19
C73 VDD sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0196f
C74 sky130_fd_sc_hd__and4_1_0/a_109_47# P2 2.77e-19
C75 G1 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0137f
C76 G4 P1 1.7e-20
C77 SUB P2 0.00318f
C78 sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/X 1.62e-19
C79 sky130_fd_sc_hd__and4_1_0/a_303_47# VDD -4.83e-19
C80 SUB sky130_fd_sc_hd__and4_1_0/X 0.251f
C81 G4 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0188f
C82 sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__a21o_1_0/X 9.17e-21
C83 SUB sky130_fd_sc_hd__a21o_1_0/X 0.461f
C84 sky130_fd_sc_hd__a21o_1_1/a_384_47# P3 7.45e-20
C85 CI P1 2.89e-19
C86 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.32e-20
C87 sky130_fd_sc_hd__and4_1_0/a_197_47# VDD -5.24e-19
C88 SUB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.0202f
C89 VDD CO -0.00363f
C90 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_1/a_384_47# 4.81e-19
C91 SUB sky130_fd_sc_hd__a21o_1_2/a_384_47# -2.27e-19
C92 SUB sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.0191f
C93 G3 SUB 6.81e-19
C94 SUB sky130_fd_sc_hd__a21o_1_3/a_81_21# -0.0199f
C95 sky130_fd_sc_hd__and4_1_0/a_109_47# P3 0.00143f
C96 VDD sky130_fd_sc_hd__a21o_1_0/a_384_47# -3.87e-19
C97 SUB P3 0.543f
C98 VDD P1 0.00652f
C99 SUB sky130_fd_sc_hd__a21o_1_2/X 0.0224f
C100 VDD sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00193f
C101 SUB P4 0.00496f
C102 sky130_fd_sc_hd__a21o_1_1/X SUB 0.0139f
C103 SUB G2 0.00126f
C104 VDD sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.0132f
C105 VDD sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00347f
C106 SUB G1 -0.00488f
C107 sky130_fd_sc_hd__and4_1_0/X P2 0.00135f
C108 SUB sky130_fd_sc_hd__a21o_1_3/a_299_297# -0.00378f
C109 SUB sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00805f
C110 sky130_fd_sc_hd__a21o_1_0/X P2 0.0752f
C111 SUB G4 8.25e-19
C112 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_0/X 7.95e-21
C113 CO P1 0.00943f
C114 P2 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00281f
C115 P2 sky130_fd_sc_hd__a21o_1_2/a_384_47# 2.47e-20
C116 sky130_fd_sc_hd__a21o_1_1/a_81_21# P2 0.0526f
C117 G3 P2 0.0287f
C118 sky130_fd_sc_hd__a21o_1_3/a_81_21# P2 6.76e-19
C119 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_2/a_384_47# 1.23e-20
C120 P1 sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.15e-20
C121 sky130_fd_sc_hd__a21o_1_3/a_81_21# sky130_fd_sc_hd__and4_1_0/X 0.0697f
C122 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.059f
C123 CI SUB 0.02f
C124 sky130_fd_sc_hd__a21o_1_1/a_384_47# VDD -4.08e-19
C125 P2 P3 0.155f
C126 SUB sky130_fd_sc_hd__a21o_1_3/a_384_47# -5.85e-20
C127 sky130_fd_sc_hd__a21o_1_2/X P2 0.455f
C128 sky130_fd_sc_hd__and4_1_0/X P3 0.00586f
C129 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_2/a_384_47# 1.12e-20
C130 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_0/X 0.0631f
C131 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__and4_1_0/X 0.132f
C132 G3 sky130_fd_sc_hd__a21o_1_0/X 0.0894f
C133 P4 P2 0.197f
C134 sky130_fd_sc_hd__a21o_1_1/X P2 0.627f
C135 P2 G2 0.00123f
C136 SUB sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00449f
C137 P4 sky130_fd_sc_hd__and4_1_0/X 4.68e-20
C138 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__and4_1_0/X 5.37e-20
C139 sky130_fd_sc_hd__a21o_1_0/X P3 0.0694f
C140 P2 G1 0.0935f
C141 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/X 0.00439f
C142 sky130_fd_sc_hd__and4_1_0/a_109_47# VDD -4.66e-19
C143 SUB sky130_fd_sc_hd__and4_1_0/a_303_47# 3.12e-20
C144 SUB VDD -0.275f
C145 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.00642f
C146 P4 sky130_fd_sc_hd__a21o_1_0/X 5.9e-20
C147 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_0/X 0.121f
C148 sky130_fd_sc_hd__and4_1_0/a_27_47# P2 0.0709f
C149 sky130_fd_sc_hd__a21o_1_0/X G2 0.0575f
C150 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/X 0.00169f
C151 G4 P2 0.00574f
C152 sky130_fd_sc_hd__a21o_1_0/X G1 0.0691f
C153 sky130_fd_sc_hd__and4_1_0/X G4 1.98e-20
C154 G3 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.023f
C155 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/a_81_21# 8.44e-20
C156 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_0/X 2.06e-20
C157 sky130_fd_sc_hd__a21o_1_2/a_384_47# P3 0.0013f
C158 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0018f
C159 sky130_fd_sc_hd__a21o_1_0/a_81_21# G2 0.0401f
C160 G3 P3 0.0176f
C161 sky130_fd_sc_hd__a21o_1_3/a_81_21# P3 2.3e-19
C162 G4 sky130_fd_sc_hd__a21o_1_0/X 3.47e-20
C163 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_2/X 0.00223f
C164 G3 sky130_fd_sc_hd__a21o_1_2/X 4.15e-19
C165 sky130_fd_sc_hd__a21o_1_3/a_81_21# sky130_fd_sc_hd__a21o_1_2/X 0.07f
C166 SUB sky130_fd_sc_hd__and4_1_0/a_197_47# -4.52e-20
C167 G1 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00416f
C168 P4 sky130_fd_sc_hd__a21o_1_2/a_384_47# 6.19e-21
C169 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_2/a_384_47# 7.94e-20
C170 SUB CO -0.00689f
C171 sky130_fd_sc_hd__a21o_1_1/a_81_21# P4 1.01e-19
C172 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0447f
C173 sky130_fd_sc_hd__a21o_1_2/X P3 0.0674f
C174 sky130_fd_sc_hd__a21o_1_1/X G3 0.0595f
C175 P4 P3 0.2f
C176 sky130_fd_sc_hd__a21o_1_1/X P3 0.185f
C177 CI P2 2.97e-20
C178 P4 sky130_fd_sc_hd__a21o_1_2/X 0.00977f
C179 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_2/X 0.0261f
C180 sky130_fd_sc_hd__a21o_1_2/X G2 5.09e-20
C181 SUB sky130_fd_sc_hd__a21o_1_0/a_384_47# -2.71e-19
C182 CI sky130_fd_sc_hd__and4_1_0/X 0.0308f
C183 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_384_47# 7.24e-19
C184 SUB P1 0.0237f
C185 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.0108f
C186 sky130_fd_sc_hd__a21o_1_1/X P4 0.0428f
C187 sky130_fd_sc_hd__a21o_1_2/X G1 4.98e-20
C188 sky130_fd_sc_hd__a21o_1_1/X G2 1.59e-19
C189 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.0173f
C190 SUB sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00449f
C191 P2 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.055f
C192 sky130_fd_sc_hd__and4_1_0/a_27_47# P3 0.0397f
C193 sky130_fd_sc_hd__a21o_1_1/X G1 0.00394f
C194 G1 G2 0.0921f
C195 SUB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.0181f
C196 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_2/X 0.0588f
C197 G4 P3 0.0694f
C198 SUB sky130_fd_sc_hd__a21o_1_0/a_299_297# -0.00449f
C199 sky130_fd_sc_hd__a21o_1_2/X G4 0.00776f
C200 sky130_fd_sc_hd__and4_1_0/a_27_47# P4 0.00576f
C201 VDD P2 0.383f
C202 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__and4_1_0/a_27_47# 1.67e-19
C203 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/X 3.17e-19
C204 SUB 0 1.71f
C205 sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C206 P1 0 0.164f
C207 P3 0 0.297f
C208 P2 0 0.31f
C209 P4 0 0.324f
C210 sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C211 CO 0 0.0276f
C212 CI 0 0.158f
C213 sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C214 sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C215 sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C216 sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C217 G4 0 0.137f
C218 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C219 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C220 sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C221 G3 0 0.137f
C222 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C223 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C224 G1 0 0.12f
C225 G2 0 0.163f
C226 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C227 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C228 VDD 0 4.61f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.25 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 A a_35_297# 0.0633f
C1 X a_35_297# 0.166f
C2 VPB a_35_297# 0.0699f
C3 a_285_297# a_35_297# 0.025f
C4 a_117_297# a_35_297# 0.00641f
C5 B a_35_297# 0.203f
C6 a_35_297# VGND 0.177f
C7 VPWR a_35_297# 0.096f
C8 X a_285_47# 0.00206f
C9 B a_285_47# 3.98e-19
C10 a_285_47# VGND 0.00552f
C11 VPWR a_285_47# 8.6e-19
C12 A X 0.00166f
C13 A VPB 0.051f
C14 VPB X 0.0154f
C15 a_35_297# a_285_47# 0.00723f
C16 A a_285_297# 0.00749f
C17 A B 0.221f
C18 a_285_297# X 0.0712f
C19 A VGND 0.0325f
C20 a_117_297# X 2.25e-19
C21 B X 0.0149f
C22 X VGND 0.173f
C23 a_285_297# VPB 0.0133f
C24 A VPWR 0.0348f
C25 B VPB 0.0697f
C26 VPB VGND 0.00696f
C27 VPWR X 0.0537f
C28 VPWR VPB 0.0689f
C29 B a_285_297# 0.0553f
C30 a_117_297# B 0.00777f
C31 a_285_297# VGND 0.00394f
C32 a_117_297# VGND 0.00177f
C33 B VGND 0.0304f
C34 a_285_297# VPWR 0.246f
C35 a_117_297# VPWR 0.00852f
C36 B VPWR 0.0703f
C37 VPWR VGND 0.0643f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt adder_3 G1 P2 G2 G3 P4 S1 S2 S3 S4 sky130_fd_sc_hd__xor2_1_3/a_117_297# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_285_47#
+ sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_117_297# CI P1 SUB
+ sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD P3
Xsky130_fd_sc_hd__xor2_1_3 P4 sky130_fd_sc_hd__xor2_1_3/B SUB SUB VDD VDD S4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a21o_1_0 CI P1 G1 SUB SUB VDD VDD sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__xor2_1_1/B P2 G2 SUB SUB VDD VDD sky130_fd_sc_hd__xor2_1_2/B
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__xor2_1_2/B P3 G3 SUB SUB VDD VDD sky130_fd_sc_hd__xor2_1_3/B
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__xor2_1_0 P1 CI SUB SUB VDD VDD S1 sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 P2 sky130_fd_sc_hd__xor2_1_1/B SUB SUB VDD VDD S2 sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 P3 sky130_fd_sc_hd__xor2_1_2/B SUB SUB VDD VDD S3 sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1
C0 S2 VDD 0.0397f
C1 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00123f
C2 sky130_fd_sc_hd__xor2_1_1/B S3 3.34e-20
C3 P1 sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.85e-19
C4 CI G2 2.73e-19
C5 SUB sky130_fd_sc_hd__a21o_1_2/a_384_47# -2.27e-19
C6 P2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0178f
C7 sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD -0.00306f
C8 S4 SUB 0.0195f
C9 CI SUB 0.176f
C10 S4 S3 0.0102f
C11 SUB P4 0.0233f
C12 S3 P4 0.00111f
C13 S1 P1 0.00593f
C14 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00109f
C15 P3 sky130_fd_sc_hd__xor2_1_1/B 0.051f
C16 G2 P2 6.94e-19
C17 S1 VDD 0.0368f
C18 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_3/B 1.77e-19
C19 SUB P2 0.384f
C20 SUB sky130_fd_sc_hd__a21o_1_0/a_384_47# 4.44e-34
C21 P3 sky130_fd_sc_hd__a21o_1_2/a_384_47# 5.7e-19
C22 sky130_fd_sc_hd__xor2_1_0/a_285_47# P1 0.00118f
C23 S1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00396f
C24 P2 S3 2.48e-20
C25 S4 P3 8.8e-19
C26 CI P3 0.346f
C27 sky130_fd_sc_hd__xor2_1_0/a_285_47# VDD -8.6e-19
C28 P3 P4 4.73e-19
C29 S2 sky130_fd_sc_hd__xor2_1_1/a_117_297# 5.82e-19
C30 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00123f
C31 G1 sky130_fd_sc_hd__xor2_1_1/B 0.0614f
C32 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0601f
C33 SUB G3 8.34e-19
C34 S2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00476f
C35 P3 P2 0.608f
C36 S4 sky130_fd_sc_hd__xor2_1_3/a_117_297# 6.67e-19
C37 sky130_fd_sc_hd__xor2_1_0/a_117_297# VDD -2.04e-19
C38 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__xor2_1_3/B 0.0322f
C39 G1 CI 0.0805f
C40 sky130_fd_sc_hd__a21o_1_0/a_299_297# P1 0.00669f
C41 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__xor2_1_2/B 0.00516f
C42 CI sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.09e-19
C43 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0562f
C44 S1 sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00102f
C45 SUB sky130_fd_sc_hd__xor2_1_2/a_35_297# -0.0113f
C46 sky130_fd_sc_hd__a21o_1_0/a_299_297# VDD 0.0016f
C47 sky130_fd_sc_hd__xor2_1_2/a_35_297# S3 0.00495f
C48 CI sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0177f
C49 S1 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0535f
C50 SUB S2 -0.00162f
C51 P2 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00611f
C52 S2 S3 0.0102f
C53 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_3/B 0.171f
C54 SUB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.0181f
C55 P3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0152f
C56 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__xor2_1_3/B 1.76e-19
C57 sky130_fd_sc_hd__xor2_1_2/a_285_297# VDD 2.35e-20
C58 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__xor2_1_2/B 4.32e-19
C59 S1 SUB -0.00328f
C60 sky130_fd_sc_hd__xor2_1_2/a_117_297# S2 8.82e-19
C61 P3 S2 0.00112f
C62 S1 S3 3.29e-19
C63 sky130_fd_sc_hd__xor2_1_1/a_285_297# S2 0.00293f
C64 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_3/B 6.06e-19
C65 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00554f
C66 P3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.57e-20
C67 SUB sky130_fd_sc_hd__xor2_1_0/a_285_47# -4.65e-19
C68 sky130_fd_sc_hd__xor2_1_0/a_285_297# VDD -3.91e-19
C69 S1 sky130_fd_sc_hd__xor2_1_2/a_117_297# 2.46e-20
C70 S1 P3 2.04e-19
C71 S1 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00137f
C72 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_384_47# 2.81e-20
C73 CI sky130_fd_sc_hd__xor2_1_1/B 0.155f
C74 SUB sky130_fd_sc_hd__xor2_1_0/a_117_297# -0.00177f
C75 sky130_fd_sc_hd__xor2_1_1/B P4 9.9e-21
C76 SUB sky130_fd_sc_hd__a21o_1_0/a_299_297# -0.00435f
C77 S4 P4 0.00239f
C78 sky130_fd_sc_hd__a21o_1_1/a_299_297# VDD 0.0016f
C79 P2 sky130_fd_sc_hd__xor2_1_1/B 0.223f
C80 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 3.85e-19
C81 SUB sky130_fd_sc_hd__xor2_1_2/a_285_297# -0.00394f
C82 sky130_fd_sc_hd__xor2_1_2/a_285_297# S3 0.00453f
C83 CI P2 0.186f
C84 CI sky130_fd_sc_hd__a21o_1_0/a_384_47# 0.00162f
C85 sky130_fd_sc_hd__xor2_1_3/B P1 0.0733f
C86 G3 sky130_fd_sc_hd__xor2_1_1/B 0.0538f
C87 sky130_fd_sc_hd__xor2_1_2/B P1 0.183f
C88 sky130_fd_sc_hd__xor2_1_3/B VDD 0.167f
C89 sky130_fd_sc_hd__xor2_1_2/B VDD 0.108f
C90 sky130_fd_sc_hd__a21o_1_1/a_384_47# VDD -4.08e-19
C91 sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00253f
C92 sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_2/B 5.8e-19
C93 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.93e-20
C94 CI G3 2.35e-19
C95 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_3/B 0.0707f
C96 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_2/B 0.00271f
C97 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_3/B 0.0593f
C98 sky130_fd_sc_hd__xor2_1_0/a_285_297# SUB -0.00394f
C99 sky130_fd_sc_hd__a21o_1_2/a_299_297# VDD 0.0344f
C100 S2 sky130_fd_sc_hd__xor2_1_1/B 0.00554f
C101 G3 P2 0.0223f
C102 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0491f
C103 sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00134f
C104 P2 sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.69e-19
C105 CI sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.2e-19
C106 S1 sky130_fd_sc_hd__xor2_1_1/B 0.112f
C107 SUB sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00436f
C108 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0714f
C109 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0151f
C110 P2 S2 0.0068f
C111 CI S1 0.002f
C112 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_0/a_285_47# 2.47e-19
C113 P2 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0197f
C114 G2 sky130_fd_sc_hd__xor2_1_3/B 2.64e-19
C115 G2 sky130_fd_sc_hd__xor2_1_2/B 0.0266f
C116 SUB sky130_fd_sc_hd__xor2_1_3/B 1.3f
C117 S1 P2 0.00354f
C118 SUB sky130_fd_sc_hd__xor2_1_2/B 0.233f
C119 sky130_fd_sc_hd__xor2_1_3/B S3 0.0617f
C120 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_1/B 0.00427f
C121 sky130_fd_sc_hd__xor2_1_2/B S3 0.00532f
C122 G3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0232f
C123 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0526f
C124 P1 VDD 0.00988f
C125 S2 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0515f
C126 P2 sky130_fd_sc_hd__xor2_1_0/a_285_47# 4.62e-19
C127 CI sky130_fd_sc_hd__xor2_1_0/a_117_297# 9.44e-19
C128 sky130_fd_sc_hd__xor2_1_0/a_35_297# P1 0.0139f
C129 S1 G3 8.29e-20
C130 sky130_fd_sc_hd__xor2_1_1/a_285_47# VDD -7.24e-19
C131 sky130_fd_sc_hd__xor2_1_2/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00134f
C132 SUB sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00449f
C133 CI sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00517f
C134 sky130_fd_sc_hd__xor2_1_2/a_117_297# sky130_fd_sc_hd__xor2_1_2/B 0.00267f
C135 P3 sky130_fd_sc_hd__xor2_1_3/B 0.159f
C136 sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 0.042f
C137 P3 sky130_fd_sc_hd__xor2_1_2/B 0.902f
C138 sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_3/B 0.00704f
C139 sky130_fd_sc_hd__xor2_1_3/a_35_297# VDD 0.00512f
C140 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_3/a_285_47# 3.65e-19
C141 S1 sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.99e-20
C142 G1 sky130_fd_sc_hd__xor2_1_3/B 1.88e-20
C143 sky130_fd_sc_hd__xor2_1_3/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00267f
C144 P3 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00623f
C145 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00303f
C146 G1 sky130_fd_sc_hd__xor2_1_2/B 0.0014f
C147 S1 S2 0.0103f
C148 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0211f
C149 sky130_fd_sc_hd__xor2_1_1/a_117_297# VDD 2.29e-20
C150 S1 sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.24e-19
C151 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.96e-19
C152 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00447f
C153 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_1/B 0.036f
C154 P1 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00101f
C155 sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00259f
C156 VDD sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00693f
C157 G2 P1 0.0104f
C158 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00128f
C159 G2 VDD 0.00129f
C160 SUB P1 1f
C161 SUB VDD -0.376f
C162 VDD S3 0.041f
C163 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__xor2_1_1/B 0.0587f
C164 SUB sky130_fd_sc_hd__xor2_1_1/a_285_47# -4.65e-19
C165 SUB sky130_fd_sc_hd__xor2_1_0/a_35_297# -0.0143f
C166 S1 sky130_fd_sc_hd__xor2_1_0/a_117_297# 4.28e-19
C167 SUB sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00517f
C168 sky130_fd_sc_hd__xor2_1_3/a_35_297# S3 0.0518f
C169 P3 P1 0.0282f
C170 S2 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00111f
C171 sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD 2.25e-20
C172 P3 VDD 0.0315f
C173 sky130_fd_sc_hd__xor2_1_3/a_285_297# S3 0.00135f
C174 sky130_fd_sc_hd__xor2_1_1/a_285_297# VDD 2.35e-20
C175 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_3/B 0.398f
C176 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_1/B 0.161f
C177 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__xor2_1_1/B 0.00123f
C178 P3 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00793f
C179 P2 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00664f
C180 SUB sky130_fd_sc_hd__xor2_1_1/a_117_297# -0.00177f
C181 sky130_fd_sc_hd__xor2_1_3/a_35_297# P3 0.00203f
C182 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__xor2_1_3/B 0.00131f
C183 sky130_fd_sc_hd__xor2_1_1/a_117_297# S3 1.88e-20
C184 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_2/a_384_47# 0.00105f
C185 S4 sky130_fd_sc_hd__xor2_1_3/B 0.00601f
C186 P1 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0152f
C187 S1 sky130_fd_sc_hd__xor2_1_2/a_285_297# 4.46e-20
C188 CI sky130_fd_sc_hd__xor2_1_3/B 0.0784f
C189 sky130_fd_sc_hd__xor2_1_3/B P4 0.104f
C190 G1 VDD 0.00163f
C191 CI sky130_fd_sc_hd__xor2_1_2/B 0.818f
C192 sky130_fd_sc_hd__xor2_1_3/a_117_297# VDD 2.25e-20
C193 VDD sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.00424f
C194 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_1/B 0.0519f
C195 SUB sky130_fd_sc_hd__xor2_1_1/a_35_297# -0.0109f
C196 P1 sky130_fd_sc_hd__a21o_1_0/a_81_21# 7.84e-20
C197 S3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 3.35e-20
C198 VDD sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00793f
C199 P2 sky130_fd_sc_hd__xor2_1_3/B 0.107f
C200 sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__xor2_1_3/B 2.82e-20
C201 P2 sky130_fd_sc_hd__xor2_1_2/B 0.163f
C202 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 1.35e-20
C203 sky130_fd_sc_hd__a21o_1_1/a_384_47# P2 6.47e-19
C204 sky130_fd_sc_hd__xor2_1_2/a_285_47# VDD -7.24e-19
C205 SUB G2 0.0237f
C206 sky130_fd_sc_hd__xor2_1_0/a_285_297# S1 0.00385f
C207 P3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.02e-19
C208 SUB S3 -0.00162f
C209 G3 sky130_fd_sc_hd__xor2_1_3/B 0.0517f
C210 G3 sky130_fd_sc_hd__xor2_1_2/B 0.0811f
C211 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_3/B 0.0908f
C212 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0262f
C213 SUB sky130_fd_sc_hd__xor2_1_2/a_117_297# -0.00177f
C214 SUB P3 0.27f
C215 sky130_fd_sc_hd__xor2_1_2/a_117_297# S3 6.67e-19
C216 P3 S3 0.00706f
C217 SUB sky130_fd_sc_hd__xor2_1_1/a_285_297# -0.00394f
C218 S1 sky130_fd_sc_hd__a21o_1_1/a_299_297# 8.32e-20
C219 sky130_fd_sc_hd__xor2_1_1/a_285_297# S3 8.64e-20
C220 S2 sky130_fd_sc_hd__xor2_1_3/B 0.0546f
C221 S2 sky130_fd_sc_hd__xor2_1_2/B 0.00962f
C222 G1 G2 1.42e-20
C223 G2 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0275f
C224 sky130_fd_sc_hd__xor2_1_1/B P1 0.132f
C225 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0563f
C226 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0116f
C227 sky130_fd_sc_hd__xor2_1_1/B VDD 0.743f
C228 G1 SUB 0.023f
C229 SUB sky130_fd_sc_hd__xor2_1_3/a_117_297# -8.18e-19
C230 SUB sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.00243f
C231 sky130_fd_sc_hd__xor2_1_3/a_117_297# S3 0.00101f
C232 G2 sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.77e-20
C233 CI P1 0.544f
C234 sky130_fd_sc_hd__a21o_1_2/a_384_47# VDD -4.08e-19
C235 S1 sky130_fd_sc_hd__xor2_1_3/B 0.0317f
C236 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_1/B 0.0678f
C237 P3 sky130_fd_sc_hd__xor2_1_3/a_285_47# 3.53e-19
C238 S1 sky130_fd_sc_hd__xor2_1_2/B 1.38e-19
C239 S4 VDD 0.0296f
C240 CI VDD 0.00219f
C241 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_1/B 5.05e-21
C242 VDD P4 0.0224f
C243 SUB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00347f
C244 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__a21o_1_2/a_384_47# 6.06e-21
C245 sky130_fd_sc_hd__xor2_1_2/a_285_47# SUB -4.65e-19
C246 CI sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0235f
C247 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00255f
C248 S4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00521f
C249 P2 P1 0.6f
C250 sky130_fd_sc_hd__a21o_1_0/a_384_47# P1 5.49e-19
C251 sky130_fd_sc_hd__xor2_1_3/a_35_297# P4 0.0132f
C252 S1 sky130_fd_sc_hd__a21o_1_2/a_299_297# 3.56e-19
C253 P2 VDD 0.0257f
C254 sky130_fd_sc_hd__a21o_1_0/a_384_47# VDD -4.08e-19
C255 S4 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.00453f
C256 sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__xor2_1_1/B 0.00269f
C257 sky130_fd_sc_hd__xor2_1_1/a_285_47# P2 0.00118f
C258 P2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00129f
C259 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/B 2.27e-19
C260 G3 P1 6.62e-19
C261 sky130_fd_sc_hd__xor2_1_2/a_285_47# P3 0.00118f
C262 sky130_fd_sc_hd__xor2_1_3/a_35_297# P2 3.67e-21
C263 G3 VDD 0.00152f
C264 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0414f
C265 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0394f
C266 G3 sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.72e-20
C267 G1 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0272f
C268 sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD 0.00796f
C269 CI sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.26e-21
C270 G2 sky130_fd_sc_hd__xor2_1_1/B 0.13f
C271 sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_3/B 0.00704f
C272 SUB sky130_fd_sc_hd__xor2_1_1/B 0.137f
C273 S3 0 0.0366f
C274 P3 0 0.733f
C275 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C276 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C277 SUB 0 1.99f
C278 S2 0 0.0353f
C279 P2 0 0.625f
C280 sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C281 VDD 0 6.64f
C282 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C283 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C284 S1 0 0.0372f
C285 P1 0 0.561f
C286 CI 0 0.811f
C287 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C288 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C289 sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C290 sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C291 G3 0 0.135f
C292 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C293 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C294 G2 0 0.134f
C295 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C296 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C297 G1 0 0.156f
C298 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C299 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C300 S4 0 0.113f
C301 P4 0 0.21f
C302 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C303 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.103 pd=0.954 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.245 ps=2.27 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.816 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.103 ps=0.954 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.136 ps=1.26 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
C0 A X 1.68e-19
C1 B VPB 0.0629f
C2 A VGND 0.0147f
C3 B X 0.00276f
C4 a_59_75# VPB 0.0563f
C5 B VGND 0.0115f
C6 a_59_75# X 0.109f
C7 X VPB 0.0127f
C8 a_59_75# VGND 0.116f
C9 a_59_75# a_145_75# 0.00658f
C10 VGND VPB 0.008f
C11 X VGND 0.0993f
C12 X a_145_75# 5.76e-19
C13 VPWR A 0.0362f
C14 VGND a_145_75# 0.00468f
C15 B VPWR 0.0117f
C16 a_59_75# VPWR 0.15f
C17 B A 0.0971f
C18 VPWR VPB 0.0729f
C19 a_59_75# A 0.0809f
C20 VPWR X 0.111f
C21 A VPB 0.0806f
C22 VPWR VGND 0.0461f
C23 a_59_75# B 0.143f
C24 VPWR a_145_75# 6.31e-19
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt adder_1 A1 B1 A2 B2 A3 B3 A4 B4 G1 P1 G2 P2 G3 P3 G4 P4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__and2_1_3/a_145_75#
+ sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__and2_1_3/a_59_75#
+ sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__and2_1_1/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__and2_1_2/a_145_75#
+ SUB sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD
Xsky130_fd_sc_hd__xor2_1_3 A4 B4 SUB SUB VDD VDD P4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 A1 B1 SUB SUB VDD VDD G1 sky130_fd_sc_hd__and2_1_0/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_1 A2 B2 SUB SUB VDD VDD G2 sky130_fd_sc_hd__and2_1_1/a_145_75#
+ sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A3 B3 SUB SUB VDD VDD G3 sky130_fd_sc_hd__and2_1_2/a_145_75#
+ sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A4 B4 SUB SUB VDD VDD G4 sky130_fd_sc_hd__and2_1_3/a_145_75#
+ sky130_fd_sc_hd__and2_1_3/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__xor2_1_0 A1 B1 SUB SUB VDD VDD P1 sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A2 B2 SUB SUB VDD VDD P2 sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A3 B3 SUB SUB VDD VDD P3 sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1
C0 VDD sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00289f
C1 A3 sky130_fd_sc_hd__xor2_1_2/a_285_297# 6.24e-19
C2 sky130_fd_sc_hd__xor2_1_2/a_35_297# A4 0.0101f
C3 A3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00595f
C4 sky130_fd_sc_hd__and2_1_0/a_59_75# A2 4.2e-20
C5 sky130_fd_sc_hd__and2_1_1/a_59_75# P1 0.00746f
C6 sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD -1.39e-19
C7 A3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 4.35e-19
C8 P1 SUB 0.0117f
C9 sky130_fd_sc_hd__and2_1_0/a_145_75# B2 1.12e-21
C10 P2 A2 0.00233f
C11 G2 VDD 0.0388f
C12 B3 A2 1e-19
C13 sky130_fd_sc_hd__and2_1_2/a_59_75# SUB 0.00617f
C14 sky130_fd_sc_hd__xor2_1_1/a_117_297# P2 5.63e-19
C15 B4 A4 0.249f
C16 sky130_fd_sc_hd__xor2_1_3/a_117_297# P4 5.63e-19
C17 P3 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.00722f
C18 P3 SUB 0.0125f
C19 G3 sky130_fd_sc_hd__and2_1_3/a_59_75# 9.08e-20
C20 VDD A2 0.198f
C21 VDD sky130_fd_sc_hd__xor2_1_3/a_117_297# -1.39e-19
C22 G2 P1 6.62e-19
C23 SUB G3 -1.95e-19
C24 P2 sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.01e-20
C25 B1 sky130_fd_sc_hd__xor2_1_0/a_285_47# 2.19e-19
C26 B4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 4.2e-19
C27 sky130_fd_sc_hd__xor2_1_3/a_35_297# P3 1.05e-19
C28 sky130_fd_sc_hd__and2_1_1/a_59_75# A3 3.22e-20
C29 sky130_fd_sc_hd__xor2_1_1/a_117_297# VDD -1.39e-19
C30 sky130_fd_sc_hd__xor2_1_3/a_35_297# G3 5.99e-22
C31 A3 SUB 0.0164f
C32 B3 G4 9.35e-20
C33 sky130_fd_sc_hd__xor2_1_2/a_117_297# P3 2.16e-19
C34 sky130_fd_sc_hd__and2_1_0/a_145_75# A1 0.00119f
C35 sky130_fd_sc_hd__xor2_1_2/a_117_297# G3 7.99e-19
C36 P1 A2 0.0305f
C37 VDD sky130_fd_sc_hd__xor2_1_0/a_285_297# 4.65e-20
C38 B2 sky130_fd_sc_hd__and2_1_1/a_145_75# 2.28e-20
C39 G2 G3 -1.94e-25
C40 P4 G4 0.00346f
C41 VDD G4 0.0395f
C42 B2 G1 7.99e-20
C43 sky130_fd_sc_hd__xor2_1_2/a_117_297# A3 0.00414f
C44 sky130_fd_sc_hd__xor2_1_1/a_117_297# P1 1.21e-19
C45 sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.6e-19
C46 G2 A3 6.19e-20
C47 sky130_fd_sc_hd__xor2_1_0/a_117_297# G1 7.26e-19
C48 sky130_fd_sc_hd__and2_1_1/a_59_75# B1 9.42e-20
C49 sky130_fd_sc_hd__xor2_1_2/a_285_297# SUB -0.00166f
C50 sky130_fd_sc_hd__xor2_1_1/a_35_297# SUB -0.00565f
C51 SUB B1 0.134f
C52 sky130_fd_sc_hd__xor2_1_3/a_117_297# P3 7.54e-20
C53 P1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00448f
C54 sky130_fd_sc_hd__xor2_1_3/a_117_297# G3 9e-22
C55 sky130_fd_sc_hd__xor2_1_3/a_285_297# G4 6.56e-19
C56 B2 A1 1.47e-19
C57 A3 A2 0.00809f
C58 sky130_fd_sc_hd__xor2_1_2/a_285_47# SUB -2.55e-19
C59 B2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 7.19e-19
C60 G2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0663f
C61 sky130_fd_sc_hd__xor2_1_0/a_117_297# A1 0.00414f
C62 G2 B1 8.95e-20
C63 G1 A1 0.0701f
C64 G2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.75e-19
C65 P3 G4 5.33e-19
C66 G1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0663f
C67 B3 A4 0.00861f
C68 G4 G3 0.00197f
C69 sky130_fd_sc_hd__and2_1_1/a_59_75# SUB 0.00649f
C70 SUB sky130_fd_sc_hd__and2_1_3/a_59_75# 0.00649f
C71 sky130_fd_sc_hd__xor2_1_1/a_35_297# A2 0.0397f
C72 sky130_fd_sc_hd__and2_1_0/a_145_75# VDD -6.31e-19
C73 A2 B1 0.00281f
C74 P4 A4 0.00232f
C75 sky130_fd_sc_hd__xor2_1_2/a_35_297# P2 1.96e-20
C76 A3 G4 1.26e-19
C77 sky130_fd_sc_hd__xor2_1_2/a_35_297# B3 0.0715f
C78 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__and2_1_3/a_59_75# 5.6e-19
C79 sky130_fd_sc_hd__xor2_1_1/a_285_297# A2 6.41e-19
C80 VDD A4 0.197f
C81 sky130_fd_sc_hd__xor2_1_3/a_35_297# SUB -0.0066f
C82 B2 sky130_fd_sc_hd__and2_1_0/a_59_75# 5.54e-20
C83 sky130_fd_sc_hd__xor2_1_0/a_35_297# A1 0.0402f
C84 sky130_fd_sc_hd__xor2_1_2/a_35_297# P4 5.81e-21
C85 sky130_fd_sc_hd__xor2_1_2/a_117_297# SUB -0.00177f
C86 sky130_fd_sc_hd__and2_1_1/a_59_75# G2 0.00228f
C87 B2 P2 0.00129f
C88 sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD 0.0079f
C89 G2 SUB -1.95e-19
C90 B2 B3 0.00271f
C91 sky130_fd_sc_hd__and2_1_0/a_59_75# G1 0.00228f
C92 sky130_fd_sc_hd__xor2_1_0/a_285_297# B1 1.19e-19
C93 sky130_fd_sc_hd__xor2_1_2/a_285_297# G4 3.71e-19
C94 B2 sky130_fd_sc_hd__xor2_1_1/a_285_47# 2.25e-19
C95 B4 B3 0.00433f
C96 sky130_fd_sc_hd__xor2_1_3/a_285_297# A4 6.41e-19
C97 sky130_fd_sc_hd__and2_1_1/a_59_75# A2 0.0589f
C98 B2 VDD 0.00698f
C99 B4 P4 0.00126f
C100 sky130_fd_sc_hd__and2_1_2/a_59_75# A4 4.2e-20
C101 A2 SUB 0.0431f
C102 sky130_fd_sc_hd__xor2_1_3/a_117_297# SUB -0.00177f
C103 VDD sky130_fd_sc_hd__and2_1_1/a_145_75# -6.31e-19
C104 sky130_fd_sc_hd__xor2_1_0/a_117_297# VDD -1.39e-19
C105 B4 VDD 0.00646f
C106 sky130_fd_sc_hd__and2_1_0/a_59_75# A1 0.0581f
C107 P3 A4 0.0296f
C108 VDD G1 0.0385f
C109 A4 G3 1.39e-19
C110 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.6e-19
C111 sky130_fd_sc_hd__xor2_1_1/a_117_297# SUB -0.00177f
C112 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__and2_1_2/a_59_75# 5.6e-19
C113 P2 A1 1.59e-21
C114 B2 P1 8.23e-19
C115 P2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.9e-21
C116 sky130_fd_sc_hd__xor2_1_2/a_35_297# P3 0.00192f
C117 A3 A4 0.00249f
C118 G2 A2 0.071f
C119 sky130_fd_sc_hd__xor2_1_2/a_35_297# G3 0.0665f
C120 sky130_fd_sc_hd__xor2_1_0/a_117_297# P1 3.4e-19
C121 sky130_fd_sc_hd__xor2_1_3/a_285_297# B4 1.19e-19
C122 G4 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0026f
C123 B2 sky130_fd_sc_hd__and2_1_2/a_59_75# 1.27e-19
C124 G4 SUB -1.95e-19
C125 P1 G1 3.4e-19
C126 VDD A1 0.182f
C127 sky130_fd_sc_hd__xor2_1_1/a_117_297# G2 7.26e-19
C128 sky130_fd_sc_hd__xor2_1_2/a_35_297# A3 0.0336f
C129 VDD sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00867f
C130 sky130_fd_sc_hd__xor2_1_3/a_35_297# G4 0.0665f
C131 B4 P3 7.42e-19
C132 G2 sky130_fd_sc_hd__xor2_1_0/a_285_297# 3.25e-19
C133 sky130_fd_sc_hd__xor2_1_2/a_285_297# A4 3.31e-19
C134 B4 G3 3.51e-20
C135 sky130_fd_sc_hd__xor2_1_2/a_117_297# G4 1.25e-19
C136 sky130_fd_sc_hd__and2_1_2/a_145_75# B2 2.37e-21
C137 B2 A3 0.00246f
C138 sky130_fd_sc_hd__xor2_1_1/a_117_297# A2 0.00414f
C139 P1 A1 0.00719f
C140 P1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00153f
C141 P2 B3 5.55e-19
C142 sky130_fd_sc_hd__xor2_1_0/a_285_297# A2 3.31e-19
C143 sky130_fd_sc_hd__and2_1_0/a_59_75# VDD -0.00241f
C144 sky130_fd_sc_hd__xor2_1_3/a_117_297# G4 7.98e-19
C145 sky130_fd_sc_hd__xor2_1_1/a_285_47# B3 3.82e-20
C146 B2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0446f
C147 B2 B1 0.00218f
C148 P2 VDD 0.0747f
C149 VDD B3 0.0264f
C150 sky130_fd_sc_hd__and2_1_3/a_145_75# A4 0.00119f
C151 B2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.19e-19
C152 B2 sky130_fd_sc_hd__xor2_1_0/a_285_47# 5.6e-20
C153 A4 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0591f
C154 A4 SUB 0.0446f
C155 G1 B1 0.0397f
C156 P1 sky130_fd_sc_hd__and2_1_0/a_59_75# 1.33e-19
C157 VDD P4 0.0238f
C158 sky130_fd_sc_hd__xor2_1_3/a_35_297# A4 0.0402f
C159 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__and2_1_3/a_59_75# 0.00179f
C160 P2 P1 3.79e-19
C161 sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB -0.0109f
C162 P2 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00164f
C163 sky130_fd_sc_hd__and2_1_1/a_59_75# B2 0.0564f
C164 A1 B1 0.264f
C165 B3 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0565f
C166 sky130_fd_sc_hd__xor2_1_3/a_285_297# P4 0.0109f
C167 B2 SUB 0.157f
C168 P1 VDD 0.0465f
C169 P2 P3 2.24e-20
C170 sky130_fd_sc_hd__and2_1_3/a_145_75# B4 2.46e-20
C171 sky130_fd_sc_hd__xor2_1_0/a_35_297# B1 0.0359f
C172 sky130_fd_sc_hd__xor2_1_3/a_285_297# VDD 2.84e-32
C173 B4 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0576f
C174 P2 G3 0.00384f
C175 P3 B3 0.00724f
C176 sky130_fd_sc_hd__xor2_1_0/a_117_297# SUB -0.00177f
C177 B4 SUB 0.154f
C178 B3 G3 0.0409f
C179 sky130_fd_sc_hd__and2_1_1/a_59_75# G1 8.11e-20
C180 sky130_fd_sc_hd__xor2_1_3/a_117_297# A4 0.00414f
C181 VDD sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00479f
C182 G1 SUB 0.00116f
C183 P2 A3 0.00732f
C184 P3 P4 2.91e-20
C185 B4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0414f
C186 A3 B3 0.294f
C187 sky130_fd_sc_hd__and2_1_2/a_145_75# B3 2.46e-20
C188 VDD P3 0.0448f
C189 B2 G2 0.042f
C190 VDD G3 0.0413f
C191 sky130_fd_sc_hd__xor2_1_0/a_117_297# G2 1.14e-19
C192 A3 P4 3.19e-21
C193 sky130_fd_sc_hd__and2_1_0/a_59_75# B1 0.0544f
C194 A3 VDD 0.208f
C195 sky130_fd_sc_hd__and2_1_2/a_145_75# VDD -6.31e-19
C196 G2 G1 0.00179f
C197 A1 SUB 0.0438f
C198 B4 sky130_fd_sc_hd__xor2_1_3/a_285_47# 2.19e-19
C199 sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00179f
C200 P2 sky130_fd_sc_hd__xor2_1_2/a_285_297# 2.5e-20
C201 P2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00234f
C202 G4 A4 0.0729f
C203 B2 A2 0.256f
C204 sky130_fd_sc_hd__xor2_1_0/a_35_297# SUB -0.00339f
C205 sky130_fd_sc_hd__xor2_1_3/a_285_297# P3 9.07e-20
C206 sky130_fd_sc_hd__xor2_1_2/a_285_297# B3 0.00523f
C207 sky130_fd_sc_hd__xor2_1_1/a_35_297# B3 4e-19
C208 P2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.0109f
C209 sky130_fd_sc_hd__and2_1_1/a_145_75# A2 0.00119f
C210 P3 sky130_fd_sc_hd__and2_1_2/a_59_75# 9.47e-20
C211 sky130_fd_sc_hd__xor2_1_2/a_285_297# P4 2.02e-20
C212 G1 A2 1.33e-19
C213 sky130_fd_sc_hd__xor2_1_2/a_35_297# G4 2.26e-19
C214 P1 A3 1.12e-21
C215 sky130_fd_sc_hd__and2_1_2/a_59_75# G3 0.0029f
C216 sky130_fd_sc_hd__xor2_1_2/a_285_297# VDD 4.65e-20
C217 VDD sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00949f
C218 G2 A1 1.14e-19
C219 VDD B1 0.00679f
C220 sky130_fd_sc_hd__xor2_1_2/a_285_47# B3 0.00257f
C221 G2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.05e-19
C222 P3 G3 2.77e-19
C223 VDD sky130_fd_sc_hd__xor2_1_1/a_285_297# 6.02e-20
C224 A3 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0594f
C225 sky130_fd_sc_hd__and2_1_0/a_59_75# SUB -0.00661f
C226 A3 P3 0.006f
C227 G1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.75e-19
C228 VDD sky130_fd_sc_hd__xor2_1_2/a_285_47# -8.2e-19
C229 B4 G4 0.0423f
C230 sky130_fd_sc_hd__and2_1_1/a_59_75# P2 4.05e-20
C231 A1 A2 0.00698f
C232 A3 G3 0.074f
C233 P1 sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.51e-19
C234 sky130_fd_sc_hd__and2_1_3/a_145_75# B3 6.15e-21
C235 P1 B1 0.0021f
C236 P2 SUB 0.00985f
C237 B3 sky130_fd_sc_hd__and2_1_3/a_59_75# 4.1e-19
C238 sky130_fd_sc_hd__xor2_1_0/a_35_297# A2 0.0101f
C239 B3 SUB 0.232f
C240 P1 sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.46e-19
C241 sky130_fd_sc_hd__and2_1_2/a_145_75# A3 0.00119f
C242 sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00133f
C243 P4 sky130_fd_sc_hd__and2_1_3/a_59_75# 2.68e-20
C244 sky130_fd_sc_hd__and2_1_3/a_145_75# VDD -6.31e-19
C245 P4 SUB 0.00985f
C246 sky130_fd_sc_hd__and2_1_1/a_59_75# VDD -7.45e-19
C247 VDD sky130_fd_sc_hd__and2_1_3/a_59_75# -7.45e-19
C248 sky130_fd_sc_hd__xor2_1_2/a_285_297# P3 0.00179f
C249 sky130_fd_sc_hd__xor2_1_1/a_35_297# P3 1.16e-20
C250 sky130_fd_sc_hd__xor2_1_2/a_117_297# P2 1.97e-20
C251 sky130_fd_sc_hd__xor2_1_0/a_285_297# A1 6.41e-19
C252 VDD SUB -0.222f
C253 sky130_fd_sc_hd__xor2_1_2/a_285_297# G3 6.58e-19
C254 G2 P2 0.00318f
C255 sky130_fd_sc_hd__xor2_1_3/a_35_297# P4 0.00234f
C256 P3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.3e-20
C257 G1 0 0.0305f
C258 SUB 0 2.81f
C259 VDD 0 7.09f
C260 P3 0 0.0173f
C261 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C262 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C263 P2 0 0.0182f
C264 A2 0 0.317f
C265 B2 0 0.338f
C266 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C267 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C268 P1 0 0.0183f
C269 A1 0 0.373f
C270 B1 0 0.337f
C271 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C272 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C273 G4 0 0.0255f
C274 B4 0 0.342f
C275 A4 0 0.328f
C276 sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C277 G3 0 0.0256f
C278 B3 0 0.339f
C279 A3 0 0.323f
C280 sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C281 G2 0 0.0255f
C282 sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C283 sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C284 P4 0 0.0763f
C285 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C286 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
.ends

.subckt adder_4 A1 B1 A2 B2 S1 S2 S3 S4 CO adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ A3 B4 adder_3_0/P4 B3 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_3_0/P3
+ adder_3_0/P2 CI adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# VDD adder_3_0/P1 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# SUB adder_2_0/G4
Xadder_2_0 CI adder_3_0/P1 adder_3_0/G1 adder_3_0/P2 adder_3_0/G2 adder_3_0/P3 adder_3_0/G3
+ adder_3_0/P4 adder_2_0/G4 CO VDD SUB adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# adder_2
Xadder_3_0 adder_3_0/G1 adder_3_0/P2 adder_3_0/G2 adder_3_0/G3 adder_3_0/P4 S1 S2
+ S3 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# CI adder_3_0/P1 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD adder_3_0/P3 adder_3
Xadder_1_0 A1 B1 A2 B2 A3 B3 A4 B4 adder_3_0/G1 adder_3_0/P1 adder_3_0/G2 adder_3_0/P2
+ adder_3_0/G3 adder_3_0/P3 adder_2_0/G4 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# SUB adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD adder_1
C0 A3 B3 1.3f
C1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B SUB -0.00596f
C2 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00465f
C3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__and4_1_0/X 6.99e-21
C4 B2 VDD 0.176f
C5 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P3 2.95e-20
C6 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -1.33e-20
C7 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/G1 6.94e-19
C8 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -2.02e-20
C9 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P1 0.00281f
C10 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G1 0.00976f
C11 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD -6.68e-19
C12 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00432f
C13 CO adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.53e-19
C14 B4 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.05e-20
C15 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P3 0.0105f
C16 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00226f
C17 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -8.72e-21
C18 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0356f
C19 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.84e-19
C20 A2 adder_3_0/G1 3.33e-19
C21 CI adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.11e-19
C22 adder_3_0/G3 B2 0.00108f
C23 adder_3_0/G2 VDD 0.293f
C24 B3 adder_2_0/G4 2.86e-19
C25 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 9.14e-21
C26 CO VDD 0.114f
C27 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# 1.86e-19
C28 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.39e-20
C29 CI VDD 1.6f
C30 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P1 1.34e-20
C31 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.11e-19
C32 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD 6.69e-20
C33 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/G3 0.00202f
C34 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.67e-19
C35 B3 A1 3.87e-19
C36 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/G1 4.07e-19
C37 adder_3_0/P2 B3 8.59e-19
C38 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# -1.01e-20
C39 adder_3_0/P4 adder_3_0/G1 1.36e-20
C40 adder_3_0/G2 adder_3_0/G3 0.882f
C41 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_2_0/G4 3.36e-19
C42 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P4 4.82e-19
C43 CO adder_3_0/G3 4.09e-20
C44 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 5.66e-20
C45 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# B3 9.41e-19
C46 CI adder_3_0/G3 0.164f
C47 A3 VDD 0.208f
C48 adder_2_0/sky130_fd_sc_hd__and4_1_0/X SUB 1.11e-19
C49 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# B3 4.89e-20
C50 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.39e-19
C51 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00611f
C52 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00131f
C53 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# adder_3_0/G1 0.00101f
C54 adder_3_0/P3 B3 0.0502f
C55 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_2_0/G4 1.03e-19
C56 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# SUB -5.32e-19
C57 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 3.54e-19
C58 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0203f
C59 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_2_0/G4 8.23e-19
C60 adder_3_0/G3 A3 0.0807f
C61 B3 adder_3_0/P1 1.06e-19
C62 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.19e-20
C63 adder_2_0/G4 VDD 0.174f
C64 A2 SUB 0.00582f
C65 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P1 0.00383f
C66 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# 8.23e-19
C67 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.14e-20
C68 A1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.52e-21
C69 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 3.36e-20
C70 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/G1 1.56e-20
C71 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# CI 0.00225f
C72 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0193f
C73 A1 VDD 0.37f
C74 B1 adder_3_0/G1 0.087f
C75 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0309f
C76 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 6.98e-20
C77 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0577f
C78 CI adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0245f
C79 adder_3_0/P2 VDD 0.267f
C80 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00125f
C81 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B S1 0.0236f
C82 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# SUB -5.69e-20
C83 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# -0.00186f
C84 adder_3_0/G3 adder_2_0/G4 0.217f
C85 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 2.22e-19
C86 adder_3_0/P4 SUB 0.492f
C87 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# VDD 0.00215f
C88 S1 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# -6.35e-20
C89 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# VDD 3.32e-19
C90 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.024f
C91 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_3_0/P3 6.88e-19
C92 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B4 3.05e-20
C93 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_2_0/G4 0.0161f
C94 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_2_0/G4 2.44e-19
C95 adder_3_0/P3 VDD 0.534f
C96 adder_3_0/G3 adder_3_0/P2 0.771f
C97 B4 A4 1.95f
C98 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/G1 3.92e-20
C99 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0275f
C100 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0208f
C101 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 5.47e-19
C102 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/G3 3.83e-19
C103 CI adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00101f
C104 adder_3_0/P1 VDD 0.332f
C105 A2 adder_3_0/P4 4.36e-19
C106 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/G3 0.0163f
C107 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.84e-20
C108 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_2_0/G4 5.98e-20
C109 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -9.51e-19
C110 adder_3_0/G3 adder_3_0/P3 0.318f
C111 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# VDD -9.12e-19
C112 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/G4 1.36e-19
C113 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00309f
C114 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_3_0/P3 0.00388f
C115 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B S2 0.118f
C116 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_3_0/P3 4.09e-20
C117 B1 SUB 0.00716f
C118 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 1.73e-19
C119 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.38e-20
C120 S1 SUB 1.38f
C121 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_3_0/G2 4.16e-19
C122 adder_2_0/sky130_fd_sc_hd__and4_1_0/X S1 0.00171f
C123 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/P2 -8.74e-21
C124 adder_3_0/G3 adder_3_0/P1 0.197f
C125 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 8.7e-19
C126 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B S4 0.0035f
C127 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0337f
C128 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B1 0.022f
C129 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/G3 -5.99e-22
C130 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 2.93e-19
C131 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.00254f
C132 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/P3 1.03e-19
C133 A2 B1 0.403f
C134 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.131f
C135 SUB adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.84e-20
C136 B4 B2 4.83e-19
C137 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD 0.00242f
C138 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00552f
C139 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00723f
C140 A1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.97e-19
C141 CI adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00104f
C142 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.39e-19
C143 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# A4 0.00264f
C144 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B4 -3.44e-20
C145 B1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00429f
C146 CI adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 2.66e-19
C147 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00437f
C148 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P1 0.0196f
C149 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# -9.88e-19
C150 S2 SUB 0.0916f
C151 adder_2_0/sky130_fd_sc_hd__and4_1_0/X S2 1.66e-20
C152 adder_3_0/P4 S1 0.00107f
C153 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0177f
C154 adder_3_0/G2 B4 9.64e-20
C155 A2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0.0155f
C156 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# adder_2_0/G4 6.97e-19
C157 B3 VDD 0.171f
C158 CI B4 1.51f
C159 S4 SUB 0.118f
C160 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# VDD 5.68e-32
C161 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00384f
C162 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -4.45e-20
C163 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/G1 0.0212f
C164 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_3_0/P2 4.8e-19
C165 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/P2 2.5e-19
C166 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.66e-20
C167 CI adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0137f
C168 A4 adder_3_0/G1 7.97e-20
C169 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 2.85e-19
C170 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/P1 0.0283f
C171 adder_3_0/G3 B3 0.0363f
C172 B4 A3 8.32e-19
C173 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00128f
C174 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B S3 0.0023f
C175 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00275f
C176 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -0.0029f
C177 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A1 9.74e-19
C178 adder_3_0/P4 S2 9.76e-19
C179 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# -9e-22
C180 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# SUB 4.59e-19
C181 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/G1 3.53e-20
C182 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X VDD 0.00147f
C183 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 2.82e-21
C184 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.82e-20
C185 B4 adder_2_0/G4 0.0886f
C186 adder_3_0/P4 S4 0.0312f
C187 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# B3 0.00199f
C188 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# -0.00268f
C189 B4 A1 2.13e-19
C190 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0105f
C191 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G1 0.017f
C192 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# -5.8e-19
C193 B4 adder_3_0/P2 9.02e-20
C194 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00197f
C195 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# SUB 9.7e-20
C196 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0407f
C197 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# SUB 1.84e-20
C198 CI adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00281f
C199 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -7.49e-19
C200 adder_3_0/G3 VDD 0.253f
C201 A4 SUB 0.00516f
C202 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# B4 3.05e-20
C203 S3 SUB 0.0886f
C204 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P2 0.00132f
C205 B2 adder_3_0/G1 2.02e-19
C206 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P1 0.00259f
C207 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# VDD -5.1e-20
C208 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.46e-20
C209 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/P1 5.17e-19
C210 B4 adder_3_0/P3 0.00132f
C211 S1 S2 1.02f
C212 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B SUB 0.00142f
C213 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.46e-21
C214 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A4 6.49e-20
C215 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.53e-19
C216 A2 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 1.08e-19
C217 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/G2 6.94e-19
C218 S1 S4 0.0283f
C219 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P3 1.5e-20
C220 B4 adder_3_0/P1 4.85e-20
C221 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# SUB 1.54e-19
C222 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -3.51e-21
C223 A2 A4 4.9e-19
C224 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_2/X -0.0153f
C225 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.34e-19
C226 adder_3_0/G2 adder_3_0/G1 0.872f
C227 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_3_0/G3 2.97e-20
C228 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# SUB -2.23e-19
C229 CI adder_3_0/G1 0.0965f
C230 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/G2 0.0946f
C231 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# CO 4.68e-19
C232 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 5.75e-20
C233 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B CO 0.477f
C234 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# B4 0.0208f
C235 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B CI -0.005f
C236 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# SUB 8.68e-19
C237 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.35e-19
C238 B2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00715f
C239 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 5.65e-19
C240 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P1 0.00658f
C241 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.00531f
C242 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B VDD -0.0577f
C243 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00591f
C244 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# SUB 4.5e-19
C245 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_2_0/G4 1.65e-19
C246 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 0.00227f
C247 adder_3_0/P4 A4 0.00541f
C248 adder_3_0/P4 S3 0.0135f
C249 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.61e-19
C250 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/G3 3.28e-19
C251 A3 adder_3_0/G1 1.32e-19
C252 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.78e-19
C253 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 6.41e-20
C254 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.92e-19
C255 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/P2 -1.11e-20
C256 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0318f
C257 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0108f
C258 B2 SUB 0.00396f
C259 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# S1 -1.76e-19
C260 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -9.62e-21
C261 S4 S2 0.0289f
C262 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB -2.36e-19
C263 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X VDD 0.0342f
C264 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# -2.26e-19
C265 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0226f
C266 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# -2.45e-19
C267 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B2 6.12e-20
C268 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00661f
C269 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.7e-20
C270 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 4.7e-20
C271 adder_3_0/G1 adder_2_0/G4 3.67e-20
C272 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/P3 0.00405f
C273 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B1 6.38e-19
C274 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.89e-20
C275 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/G4 8.62e-20
C276 adder_3_0/G2 SUB 0.287f
C277 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.49e-19
C278 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# A3 9.09e-19
C279 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0.106f
C280 CO SUB 0.151f
C281 A2 B2 0.77f
C282 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/P2 0.00105f
C283 CI SUB 1.48f
C284 CI adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0.0231f
C285 adder_3_0/G1 A1 0.0955f
C286 B1 A4 3.49e-19
C287 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.71e-20
C288 SUB adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 4.55e-19
C289 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00133f
C290 adder_3_0/P2 adder_3_0/G1 0.268f
C291 S3 S1 0.0279f
C292 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P2 -0.0409f
C293 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 5.12e-19
C294 B4 B3 8.66e-19
C295 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G2 0.00105f
C296 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 4.64e-20
C297 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00898f
C298 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0151f
C299 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 7.13e-21
C300 A2 adder_3_0/G2 0.084f
C301 adder_3_0/P4 B2 6.88e-19
C302 adder_2_0/sky130_fd_sc_hd__and4_1_0/X A3 3.53e-20
C303 A3 SUB 0.00693f
C304 adder_3_0/P3 adder_3_0/G1 8.5e-20
C305 A2 CI 2.43e-19
C306 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# adder_3_0/P3 4.99e-19
C307 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P3 0.00276f
C308 S1 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 9.19e-19
C309 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.92e-20
C310 S1 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 6.31e-20
C311 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 0.00366f
C312 A4 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.72e-20
C313 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# S3 9.42e-19
C314 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00176f
C315 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A3 1e-19
C316 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/P2 0.0124f
C317 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# SUB 7.61e-19
C318 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/G2 7.19e-20
C319 adder_3_0/G1 adder_3_0/P1 0.0488f
C320 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# S1 -0.00115f
C321 CI adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.0208f
C322 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# adder_3_0/P1 2.07e-19
C323 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 0.00637f
C324 adder_3_0/P4 adder_3_0/G2 4.99e-20
C325 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P1 0.103f
C326 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00297f
C327 CO adder_3_0/P4 6.01e-19
C328 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_2_0/G4 1.36e-19
C329 A2 A3 0.00214f
C330 SUB adder_2_0/G4 0.132f
C331 adder_3_0/P4 CI 0.0664f
C332 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 4.86e-19
C333 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S4 0.00104f
C334 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/G1 0.0118f
C335 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P1 1.85e-21
C336 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P2 1.63e-19
C337 S3 S2 0.717f
C338 S1 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -2.34e-19
C339 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# 5.09e-21
C340 SUB A1 0.00365f
C341 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.27e-21
C342 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 2.6e-21
C343 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/P4 0.00212f
C344 adder_3_0/P2 SUB 0.0707f
C345 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# S4 -3.24e-19
C346 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P2 -2.14e-20
C347 B1 B2 0.00145f
C348 B4 VDD 0.138f
C349 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0283f
C350 S3 S4 0.442f
C351 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.84e-32
C352 adder_3_0/P4 A3 1.54e-19
C353 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# SUB 1.4e-19
C354 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A1 -6.08e-19
C355 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 7.89e-20
C356 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P3 0.0039f
C357 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/P1 3.68e-21
C358 A2 adder_2_0/G4 1.33e-19
C359 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.00146f
C360 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# SUB 3.52e-21
C361 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_2_0/sky130_fd_sc_hd__and4_1_0/X 7.41e-22
C362 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P2 2.17e-19
C363 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 7.63e-20
C364 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P3 5.85e-19
C365 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# B3 0.0195f
C366 adder_3_0/P3 SUB 0.136f
C367 A2 A1 0.00288f
C368 B4 adder_3_0/G3 9.64e-20
C369 B1 adder_3_0/G2 0.00409f
C370 CI adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 1.5e-20
C371 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/P4 4.5e-19
C372 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.44e-19
C373 A2 adder_3_0/P2 0.00581f
C374 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# S2 0.00567f
C375 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P1 5.1e-19
C376 CI B1 1.95e-19
C377 CO S1 0.257f
C378 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.0072f
C379 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# B4 5.56e-19
C380 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# S2 9.42e-19
C381 CI S1 4.68e-19
C382 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.77e-19
C383 B2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 6.16e-19
C384 adder_3_0/P4 adder_2_0/G4 1.29f
C385 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# -7.29e-19
C386 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P1 0.00468f
C387 SUB adder_3_0/P1 0.175f
C388 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P3 5.23e-19
C389 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# SUB 8.85e-19
C390 A2 adder_3_0/P3 2.27e-19
C391 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# S1 -3.09e-20
C392 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# SUB 9.8e-19
C393 adder_3_0/P4 adder_3_0/P2 0.0172f
C394 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/P1 0.00105f
C395 B1 A3 9.01e-19
C396 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P1 0.0152f
C397 B3 adder_3_0/G1 1.01e-19
C398 CI adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# 9.49e-19
C399 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0.0173f
C400 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB 6.56e-19
C401 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/G1 3.22e-19
C402 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.55e-19
C403 CI adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.01e-20
C404 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.04e-19
C405 A2 adder_3_0/P1 0.0449f
C406 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.55e-20
C407 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A4 3.72e-20
C408 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S3 7.3e-19
C409 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 9.82e-21
C410 adder_3_0/P4 adder_3_0/P3 0.232f
C411 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# S1 -1.39e-20
C412 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.99e-19
C413 CO S2 0.0426f
C414 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_3_0/P1 0.00143f
C415 CI S2 0.00387f
C416 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/P1 3.41e-19
C417 S1 adder_2_0/G4 2.86e-20
C418 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 3.33e-20
C419 A3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 5.96e-20
C420 adder_3_0/P4 adder_3_0/P1 0.0308f
C421 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.04e-19
C422 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.0141f
C423 B1 A1 0.237f
C424 CO S4 0.209f
C425 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.045f
C426 B1 adder_3_0/P2 6.78e-19
C427 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/G3 2.64e-19
C428 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/P4 0.0131f
C429 S1 adder_3_0/P2 0.234f
C430 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 2.56e-19
C431 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 1.03e-19
C432 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A4 6.49e-20
C433 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00475f
C434 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# S1 1.21e-20
C435 adder_3_0/G1 VDD 0.694f
C436 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# -4.4e-19
C437 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00101f
C438 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/G4 1.82e-19
C439 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B VDD -0.019f
C440 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 8.63e-21
C441 adder_2_0/sky130_fd_sc_hd__and4_1_0/X B3 1.55e-20
C442 SUB B3 0.00596f
C443 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 9.74e-19
C444 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 6.84e-21
C445 S1 adder_3_0/P3 0.1f
C446 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.21e-19
C447 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 5.64e-19
C448 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X -1.77e-19
C449 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B3 7.98e-20
C450 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/G2 1.77e-21
C451 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B2 7.88e-20
C452 B1 adder_3_0/P1 0.0278f
C453 adder_3_0/G3 adder_3_0/G1 0.0163f
C454 S2 adder_2_0/G4 2.28e-20
C455 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.5e-20
C456 CI adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.49e-19
C457 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 3.35e-21
C458 S1 adder_3_0/P1 0.0451f
C459 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# -4.62e-19
C460 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/G3 0.00104f
C461 B2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00385f
C462 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.73e-19
C463 B2 A4 8.41e-19
C464 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# 3.18e-19
C465 CI adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# 3.82e-20
C466 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.13e-20
C467 A2 B3 7.94e-19
C468 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_3_0/P3 9.41e-19
C469 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# VDD 5.68e-32
C470 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 4.76e-20
C471 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00352f
C472 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_3_0/P3 1.14e-19
C473 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 5.59e-20
C474 S2 adder_3_0/P2 0.0771f
C475 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A4 0.00128f
C476 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00249f
C477 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/G4 0.00559f
C478 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G2 0.0185f
C479 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/G2 7.89e-19
C480 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S1 3.79e-19
C481 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# VDD -5.68e-32
C482 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CI 2.96e-20
C483 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# B3 4.93e-21
C484 CI adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.82e-19
C485 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 4.07e-19
C486 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -6.74e-19
C487 adder_3_0/G2 A4 1.16e-19
C488 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00285f
C489 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/P1 0.00384f
C490 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.82e-20
C491 adder_3_0/P4 B3 1.46e-19
C492 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# B2 5.71e-20
C493 adder_3_0/P3 S2 0.238f
C494 B2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.92e-20
C495 CI A4 0.0346f
C496 adder_2_0/sky130_fd_sc_hd__and4_1_0/X VDD -0.0032f
C497 SUB VDD 1.2f
C498 CO S3 0.119f
C499 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B2 0.0195f
C500 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0407f
C501 S4 adder_3_0/P3 -8.8e-19
C502 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 5.31e-21
C503 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -0.014f
C504 CO adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0228f
C505 CI adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.31e-19
C506 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A3 5.96e-20
C507 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD -4.41e-19
C508 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/G4 0.00122f
C509 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 9.54e-19
C510 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/P3 0.00147f
C511 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 1.47e-20
C512 A3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 2.11e-19
C513 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 4.68e-20
C514 adder_3_0/G3 SUB 1.22f
C515 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.74e-19
C516 A3 A4 0.00106f
C517 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00806f
C518 CI adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00244f
C519 CO adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0284f
C520 CI adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0104f
C521 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00912f
C522 A2 VDD 0.227f
C523 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S4 -1.86e-19
C524 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 1.69e-19
C525 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.45e-19
C526 CI adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.53e-20
C527 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# SUB 3.16e-20
C528 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P2 0.00106f
C529 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00776f
C530 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.014f
C531 CI adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00503f
C532 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# 0.00103f
C533 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S2 0.00273f
C534 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G3 0.00129f
C535 B1 B3 5.26e-19
C536 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0445f
C537 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G2 0.00133f
C538 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00539f
C539 B1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00727f
C540 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 1.8e-19
C541 CI adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0052f
C542 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 6.98e-20
C543 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 4e-19
C544 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 3.05e-20
C545 A2 adder_3_0/G3 0.0115f
C546 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_2_0/G4 3.67e-19
C547 A4 adder_2_0/G4 0.0821f
C548 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A1 0.0155f
C549 A3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 5.54e-20
C550 adder_3_0/P4 VDD 0.896f
C551 CO adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 1.62e-20
C552 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A1 0.00131f
C553 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P3 0.00509f
C554 S3 adder_2_0/G4 2.78e-20
C555 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.6e-20
C556 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A3 5.49e-19
C557 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P2 -1.88e-20
C558 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# adder_3_0/P3 4.98e-19
C559 A4 A1 2.8e-19
C560 adder_3_0/G2 B2 0.089f
C561 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/G4 0.00256f
C562 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# VDD 8.07e-19
C563 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00103f
C564 CI B2 3.41e-19
C565 A4 adder_3_0/P2 1.08e-19
C566 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# 8.25e-19
C567 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.00204f
C568 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 7.03e-19
C569 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00238f
C570 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 3.12e-19
C571 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# B3 5.14e-19
C572 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P1 2.37e-21
C573 S3 adder_3_0/P2 3.05e-21
C574 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 9.34e-21
C575 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/G2 1.11e-21
C576 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# -2.17e-19
C577 adder_3_0/P4 adder_3_0/G3 0.00126f
C578 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# B3 4.65e-20
C579 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# adder_3_0/P3 -3.53e-19
C580 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# CI 0.0185f
C581 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_2_0/G4 1.75e-19
C582 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P3 5.91e-19
C583 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_2_0/G4 0.0203f
C584 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.00628f
C585 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# A4 3.72e-20
C586 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/G4 7.97e-20
C587 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.011f
C588 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 4.95e-20
C589 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.99e-19
C590 adder_3_0/P3 A4 0.0462f
C591 B2 A3 0.938f
C592 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/G4 1.23e-20
C593 CI adder_3_0/G2 0.0259f
C594 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.37e-21
C595 S3 adder_3_0/P3 0.0899f
C596 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 3.97e-19
C597 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P2 4.11e-19
C598 CO CI 0.0904f
C599 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0146f
C600 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0208f
C601 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00441f
C602 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/P1 -6e-21
C603 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P1 0.00383f
C604 CI adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00313f
C605 B1 VDD 0.244f
C606 CI adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.49e-19
C607 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P2 0.0148f
C608 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A3 -7.46e-20
C609 S1 VDD -0.00292f
C610 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -0.00685f
C611 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 6.92e-20
C612 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/P1 3.02e-21
C613 A4 adder_3_0/P1 8.78e-20
C614 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 9.53e-20
C615 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G1 0.0239f
C616 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# CO 6.62e-19
C617 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 6.41e-20
C618 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 8.48e-19
C619 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# -7.21e-19
C620 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/G1 4.44e-19
C621 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.09e-19
C622 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P3 0.00835f
C623 adder_3_0/G2 A3 2.08e-19
C624 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# A4 -2.86e-19
C625 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.05e-20
C626 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0225f
C627 B2 adder_2_0/G4 0.00161f
C628 CO A3 0.00124f
C629 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P1 -6.47e-19
C630 CI A3 0.0954f
C631 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.5e-19
C632 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 8.3e-19
C633 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P3 0.00106f
C634 B1 adder_3_0/G3 0.00439f
C635 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0026f
C636 adder_3_0/G3 S1 6.53e-19
C637 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 4.59e-19
C638 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# VDD -8.51e-21
C639 B4 adder_3_0/G1 6.45e-20
C640 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P3 1.78e-19
C641 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# CO 3.28e-19
C642 B2 A1 9.29e-19
C643 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# CI 6.1e-19
C644 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_2_0/G4 1.9e-19
C645 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P1 0.0174f
C646 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# VDD 2.99e-19
C647 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S3 0.00559f
C648 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/P1 0.0274f
C649 B2 adder_3_0/P2 0.0325f
C650 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P3 5.63e-21
C651 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# CO 4.34e-19
C652 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00229f
C653 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.81e-19
C654 CI adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.33e-19
C655 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P1 1.38e-19
C656 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0383f
C657 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -0.00152f
C658 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/G1 0.00311f
C659 adder_3_0/G2 adder_2_0/G4 7.19e-19
C660 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P1 -9.58e-19
C661 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P2 -9.82e-21
C662 CO adder_2_0/G4 1.56e-19
C663 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# -0.00512f
C664 CI adder_2_0/G4 0.0329f
C665 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0084f
C666 S2 VDD 0.00253f
C667 adder_3_0/G2 A1 0.00324f
C668 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P1 7.78e-20
C669 B2 adder_3_0/P3 0.00568f
C670 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0.00261f
C671 CI A1 1.72e-19
C672 adder_3_0/G2 adder_3_0/P2 0.749f
C673 CO adder_3_0/P2 0.108f
C674 CI adder_3_0/P2 0.0316f
C675 S4 VDD -2.22e-19
C676 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P3 0.011f
C677 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00225f
C678 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 9.07e-20
C679 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.00968f
C680 B2 adder_3_0/P1 0.00166f
C681 A3 adder_2_0/G4 2.73e-19
C682 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 7.55e-22
C683 CO adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00874f
C684 CI adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.0104f
C685 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/G2 1.78e-20
C686 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00216f
C687 CO adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.8e-20
C688 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B3 4.65e-20
C689 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# 6.85e-19
C690 CI adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 5.48e-19
C691 adder_3_0/G2 adder_3_0/P3 0.0027f
C692 A3 A1 5.77e-19
C693 CO adder_3_0/P3 0.0888f
C694 CI adder_3_0/P3 0.132f
C695 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 0.00104f
C696 A4 B3 1.7f
C697 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/P3 1.36e-19
C698 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.7e-19
C699 A3 adder_3_0/P2 0.0346f
C700 B4 SUB 0.00678f
C701 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/G4 1.01e-20
C702 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# adder_3_0/P2 4.99e-19
C703 adder_3_0/G2 adder_3_0/P1 0.405f
C704 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A3 2.34e-21
C705 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/P3 3.13e-19
C706 CO adder_3_0/P1 0.0294f
C707 CI adder_3_0/P1 0.154f
C708 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 9.58e-21
C709 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.31e-20
C710 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# A3 0.0163f
C711 adder_3_0/P1 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 5.85e-19
C712 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B4 5.38e-20
C713 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P2 -8.11e-19
C714 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD 1.34e-19
C715 adder_3_0/P3 A3 0.002f
C716 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/G2 0.0051f
C717 CI adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 4.51e-20
C718 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X B3 1.6e-20
C719 adder_3_0/P2 adder_2_0/G4 0.0231f
C720 A2 B4 3.27e-19
C721 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B3 2.25e-20
C722 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0038f
C723 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 7.73e-19
C724 adder_3_0/P2 A1 3.75e-19
C725 B2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 8.1e-20
C726 A3 adder_3_0/P1 1.31e-19
C727 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_2_0/G4 1.75e-19
C728 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P3 0.00801f
C729 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -4.9e-21
C730 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_2_0/G4 4.89e-20
C731 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00612f
C732 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/G3 0.0147f
C733 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# VDD 0.00935f
C734 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD 0.00221f
C735 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 7.32e-20
C736 adder_3_0/P3 adder_2_0/G4 1.15f
C737 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P2 0.00114f
C738 adder_3_0/P4 B4 0.0321f
C739 A4 VDD 0.142f
C740 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P1 7.47e-19
C741 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/G1 -6.76e-19
C742 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/P2 0.00223f
C743 S3 VDD 8.27e-19
C744 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 9.85e-20
C745 adder_3_0/P3 adder_3_0/P2 0.405f
C746 B2 B3 0.00119f
C747 adder_3_0/P1 adder_2_0/G4 0.03f
C748 CI adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.83e-19
C749 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B VDD -2.88e-19
C750 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 1.13e-19
C751 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G3 0.00395f
C752 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00349f
C753 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P3 1.34e-19
C754 A1 adder_3_0/P1 0.00472f
C755 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 8.67e-21
C756 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B3 0.0107f
C757 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.69e-19
C758 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_2_0/G4 0.00895f
C759 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# SUB -5.95e-20
C760 adder_3_0/G3 A4 1.67e-19
C761 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 8.1e-20
C762 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/P3 7.39e-20
C763 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# VDD 0.00235f
C764 adder_3_0/P2 adder_3_0/P1 1.17f
C765 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X VDD 0.00224f
C766 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD -6.01e-19
C767 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# A4 0.0161f
C768 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -8.36e-21
C769 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_2_0/G4 3.23e-20
C770 adder_3_0/G2 B3 1.49e-19
C771 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0127f
C772 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P1 0.00112f
C773 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD 4.68e-19
C774 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P2 0.00724f
C775 CI B3 0.208f
C776 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.95e-19
C777 B1 B4 2.5e-19
C778 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 6.51e-19
C779 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.99e-20
C780 adder_3_0/P3 adder_3_0/P1 0.649f
C781 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 3.99e-20
C782 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P2 -4.84e-19
C783 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0333f
C784 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# VDD -0.00753f
C785 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/G3 4.15e-19
C786 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P2 0.00242f
C787 SUB adder_3_0/G1 0.376f
C788 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/P3 3.07e-20
C789 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 3.16e-19
C790 B2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.07e-20
C791 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C792 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C793 A2 0 0.553f
C794 B2 0 0.632f
C795 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C796 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C797 A1 0 0.469f
C798 B1 0 0.496f
C799 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C800 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C801 B4 0 1.05f
C802 A4 0 0.714f
C803 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C804 B3 0 0.683f
C805 A3 0 0.729f
C806 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C807 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C808 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C809 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C810 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C811 S3 0 0.233f
C812 adder_3_0/P3 0 1.49f
C813 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C814 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C815 SUB 0 8.51f
C816 S2 0 0.212f
C817 adder_3_0/P2 0 1.26f
C818 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C819 VDD 0 17.6f
C820 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C821 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C822 S1 0 0.285f
C823 adder_3_0/P1 0 1.11f
C824 CI 0 2.13f
C825 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C826 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C827 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C828 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C829 adder_3_0/G3 0 0.718f
C830 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C831 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C832 adder_3_0/G2 0 0.642f
C833 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C834 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C835 adder_3_0/G1 0 0.527f
C836 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C837 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C838 S4 0 0.335f
C839 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C840 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C841 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C842 adder_3_0/P4 0 1.62f
C843 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C844 CO 0 0.959f
C845 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C846 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C847 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C848 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C849 adder_2_0/G4 0 0.596f
C850 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C851 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C852 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C853 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C854 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C855 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C856 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

.subckt adder A1 B1 A2 B2 A3 B3 A4 B4 A5 B5 A6 B6 A7 B7 A8 B8 A9 B9 A10 B10 A11 B11
+ A12 B12 A13 B13 A14 B14 A15 B15 A16 B16 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13
+ S14 S15 S16 CI CO VDD GND
Xadder_4_1 A5 B5 A6 B6 S5 S6 S7 S8 adder_4_2/CI adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_1/adder_3_0/G3
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_1/adder_3_0/G2
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_1/adder_3_0/G1 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A8 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ A7 B8 adder_4_1/adder_3_0/P4 B7 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75#
+ adder_4_1/adder_3_0/P3 adder_4_1/adder_3_0/P2 adder_4_1/CI adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ VDD adder_4_1/adder_3_0/P1 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND adder_4_1/adder_2_0/G4
+ adder_4
Xadder_4_2 A9 B9 A10 B10 S9 S10 S11 S12 adder_4_3/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_2/adder_3_0/G3
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_2/adder_3_0/G2
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_2/adder_3_0/G1 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A12 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ A11 B12 adder_4_2/adder_3_0/P4 B11 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75#
+ adder_4_2/adder_3_0/P3 adder_4_2/adder_3_0/P2 adder_4_2/CI adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ VDD adder_4_2/adder_3_0/P1 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND adder_4_2/adder_2_0/G4
+ adder_4
Xadder_4_3 A13 B13 A14 B14 S13 S14 S15 S16 CO adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_3/adder_3_0/G3
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_3/adder_3_0/G2
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/adder_3_0/G1 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A16 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ A15 B16 adder_4_3/adder_3_0/P4 B15 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75#
+ adder_4_3/adder_3_0/P3 adder_4_3/adder_3_0/P2 adder_4_3/CI adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ VDD adder_4_3/adder_3_0/P1 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND adder_4_3/adder_2_0/G4
+ adder_4
Xadder_4_0 A1 B1 A2 B2 S1 S2 S3 S4 adder_4_1/CI adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_0/adder_3_0/G3
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_0/adder_3_0/G2
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_0/adder_3_0/G1 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A4 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ A3 B4 adder_4_0/adder_3_0/P4 B3 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75#
+ adder_4_0/adder_3_0/P3 adder_4_0/adder_3_0/P2 CI adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ VDD adder_4_0/adder_3_0/P1 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND adder_4_0/adder_2_0/G4
+ adder_4
C0 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# A12 6.43e-20
C1 A8 VDD 0.0408f
C2 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.74e-19
C3 S8 GND 6.99e-20
C4 B5 adder_4_0/adder_3_0/P1 8.38e-20
C5 A14 adder_4_2/adder_3_0/P1 1.27e-19
C6 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.64e-20
C7 A8 GND 0.00203f
C8 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.28e-21
C9 B16 S11 4.77e-19
C10 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.433f
C11 adder_4_0/adder_3_0/G3 VDD 5.85e-20
C12 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B16 1.66e-19
C13 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B5 1.56e-20
C14 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.46e-19
C15 B11 adder_4_1/adder_3_0/G1 9.39e-20
C16 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.7e-20
C17 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00191f
C18 GND adder_4_0/adder_3_0/G3 -1.42e-32
C19 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A12 1.39e-19
C20 B16 adder_4_2/CI 7.74e-19
C21 adder_4_1/CI adder_4_2/adder_3_0/P1 2.44e-20
C22 B11 adder_4_1/adder_3_0/P3 2.06e-19
C23 A6 adder_4_0/adder_3_0/G3 8.92e-19
C24 A9 VDD 0.0675f
C25 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.42e-19
C26 adder_4_1/adder_3_0/P3 adder_4_2/adder_3_0/G3 2.38e-20
C27 CI A7 2.75e-19
C28 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# VDD 4.75e-20
C29 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C30 B8 adder_4_0/adder_3_0/P2 4.43e-19
C31 adder_4_2/adder_3_0/P2 B14 1.84e-19
C32 A9 GND 1.99e-19
C33 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 8.75e-20
C34 S1 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.99e-21
C35 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.39e-19
C36 adder_4_2/adder_3_0/P2 B15 3.03e-19
C37 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.8e-21
C38 adder_4_0/adder_3_0/P1 A5 2.83e-20
C39 adder_4_3/CI adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 4.64e-20
C40 B7 VDD 0.0408f
C41 adder_4_2/adder_3_0/P2 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.18e-20
C42 adder_4_1/adder_3_0/P2 adder_4_0/adder_3_0/P3 2.36e-20
C43 B8 adder_4_0/adder_3_0/G1 1.31e-19
C44 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.19e-20
C45 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A5 2.25e-19
C46 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.8e-20
C47 B7 GND 0.00112f
C48 adder_4_2/adder_3_0/P2 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.19e-20
C49 S9 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.99e-21
C50 adder_4_3/adder_3_0/P1 adder_4_2/adder_3_0/P2 0.00296f
C51 adder_4_1/adder_3_0/P3 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.97e-20
C52 adder_4_1/CI A10 1.92e-19
C53 A16 S10 1.69e-19
C54 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# VDD 4.75e-20
C55 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/P2 2.08e-20
C56 adder_4_2/adder_3_0/P3 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.44e-19
C57 adder_4_2/adder_2_0/G4 GND 4.83e-20
C58 adder_4_3/CI adder_4_2/adder_3_0/G3 1.54e-19
C59 S1 A8 1.3e-19
C60 adder_4_2/adder_3_0/P2 adder_4_3/adder_3_0/G2 6.64e-21
C61 CI adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.8e-20
C62 A15 adder_4_2/adder_3_0/P3 2.29e-19
C63 adder_4_0/adder_3_0/P1 B6 1.48e-19
C64 A8 S4 3.33e-19
C65 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# CI 2.46e-19
C66 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 5.65e-20
C67 S5 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.99e-21
C68 adder_4_1/adder_2_0/G4 S3 2.25e-20
C69 A12 VDD 0.0408f
C70 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 7.91e-21
C71 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B6 2.01e-20
C72 S9 B15 8.93e-20
C73 adder_4_0/adder_3_0/G2 B8 1.21e-19
C74 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.18e-19
C75 adder_4_1/CI CI 0.0496f
C76 GND adder_4_3/adder_3_0/G3 5.02e-20
C77 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# GND 7.65e-19
C78 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.39e-35
C79 GND A12 0.00154f
C80 adder_4_1/CI adder_4_1/adder_3_0/P3 3.24e-20
C81 A7 adder_4_0/adder_3_0/P2 1.97e-19
C82 adder_4_1/adder_3_0/G1 A10 6.2e-20
C83 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.76e-20
C84 adder_4_2/adder_3_0/G1 B16 1.31e-19
C85 adder_4_1/adder_2_0/G4 adder_4_2/CI 1.64e-21
C86 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.72e-21
C87 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A12 4.77e-20
C88 A10 adder_4_1/adder_3_0/P3 4.46e-20
C89 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S11 2.47e-20
C90 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.2e-20
C91 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.78e-20
C92 adder_4_3/CI adder_4_2/adder_3_0/P1 4.71e-19
C93 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 5e-21
C94 adder_4_0/adder_3_0/G1 A7 8.1e-20
C95 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A8 3.71e-19
C96 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B14 2.06e-22
C97 adder_4_1/adder_3_0/G2 B9 1.61e-19
C98 B8 adder_4_0/adder_3_0/P3 5.72e-19
C99 S11 adder_4_3/adder_3_0/P4 2.35e-20
C100 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.32e-20
C101 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B15 4.06e-20
C102 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 2.02e-19
C103 S1 B7 8.93e-20
C104 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00977f
C105 adder_4_3/adder_3_0/P3 S9 1.67e-20
C106 A5 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.68e-19
C107 adder_4_3/adder_3_0/G1 adder_4_2/adder_3_0/P1 7.91e-22
C108 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.29e-19
C109 adder_4_2/adder_3_0/P4 S8 2.69e-20
C110 adder_4_1/adder_3_0/P1 VDD 0.00153f
C111 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_4_3/CI 2.13e-21
C112 B8 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.93e-22
C113 adder_4_2/adder_3_0/G3 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.18e-20
C114 CI adder_4_1/adder_3_0/G1 0.0031f
C115 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_4_2/CI 4.91e-21
C116 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# GND 1.66e-20
C117 adder_4_0/adder_3_0/P2 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.6e-19
C118 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S7 5.56e-20
C119 B5 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00399f
C120 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S6 1.18e-20
C121 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD 4.95e-20
C122 A11 adder_4_1/adder_3_0/P1 1.89e-19
C123 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.79e-20
C124 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B VDD 1.37e-19
C125 adder_4_0/adder_3_0/G2 A7 7.47e-20
C126 A1 VDD 1.39e-19
C127 adder_4_2/adder_3_0/G2 VDD 4.62e-20
C128 adder_4_1/CI adder_4_0/adder_3_0/P2 6.08e-19
C129 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD 4.95e-20
C130 S12 B16 5.46e-19
C131 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B7 2.9e-20
C132 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# S11 1.39e-20
C133 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.01e-20
C134 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.14e-19
C135 S1 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.6e-21
C136 adder_4_2/adder_3_0/G2 GND 1.6e-20
C137 S3 VDD 2.72e-19
C138 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# GND 1.01e-20
C139 adder_4_1/CI adder_4_0/adder_3_0/G1 1.58e-19
C140 adder_4_1/adder_2_0/G4 B12 1.47e-21
C141 B8 S2 3.18e-19
C142 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S4 7.81e-20
C143 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_2/adder_3_0/P1 2.81e-20
C144 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 3.81e-20
C145 S11 VDD 2.72e-19
C146 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B VDD 0.0303f
C147 B10 VDD 0.0407f
C148 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.28e-21
C149 GND S3 0.0398f
C150 A7 adder_4_0/adder_3_0/P3 2.29e-19
C151 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.66e-19
C152 A5 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.79e-20
C153 B10 GND 6.79e-19
C154 adder_4_2/CI VDD 0.156f
C155 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B A10 1.53e-19
C156 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_1/adder_3_0/G3 2.84e-32
C157 CI adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.01e-20
C158 adder_4_2/CI GND 0.04f
C159 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B10 2.06e-22
C160 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.43e-20
C161 B13 VDD 0.0449f
C162 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# GND 1.76e-20
C163 B7 adder_4_1/adder_3_0/G2 1.39e-35
C164 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 9.13e-20
C165 B16 adder_4_2/adder_3_0/G3 1.27e-19
C166 S5 adder_4_2/adder_2_0/G4 1.75e-20
C167 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X B12 4.4e-21
C168 A11 adder_4_2/CI 0.00338f
C169 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_2/CI 6.87e-20
C170 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# GND 1.39e-20
C171 S1 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 5.99e-21
C172 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.29e-19
C173 GND B13 1.84e-19
C174 adder_4_2/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 2.86e-20
C175 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# GND 1.39e-20
C176 adder_4_1/CI adder_4_0/adder_3_0/G2 1.47e-19
C177 B14 VDD 0.0407f
C178 A13 VDD 0.0675f
C179 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# GND 1.99e-19
C180 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.01e-20
C181 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.05e-19
C182 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S10 5.48e-20
C183 B15 VDD 0.0408f
C184 GND B14 6.79e-19
C185 B5 CI 1.09e-19
C186 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.32e-20
C187 A13 GND 1.99e-19
C188 adder_4_3/adder_3_0/P2 adder_4_2/CI 4.97e-20
C189 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_2/adder_3_0/P1 2.06e-19
C190 S2 adder_4_1/adder_3_0/P4 2.06e-20
C191 S2 A7 3.71e-20
C192 B15 GND 0.00112f
C193 S5 A12 1.3e-19
C194 A14 adder_4_2/adder_3_0/P2 1.62e-19
C195 A15 S10 3.71e-20
C196 adder_4_1/adder_2_0/G4 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 9.08e-21
C197 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# GND 1.39e-20
C198 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/CI 0.433f
C199 adder_4_1/CI adder_4_0/adder_3_0/P3 7.78e-19
C200 B16 adder_4_2/adder_3_0/P1 3.59e-19
C201 adder_4_1/adder_3_0/G2 A12 1.02e-19
C202 adder_4_1/adder_3_0/P2 VDD 9.04e-19
C203 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND 1.39e-20
C204 B8 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.4e-21
C205 adder_4_3/adder_2_0/G4 adder_4_3/CI 3.53e-20
C206 adder_4_0/adder_3_0/P1 VDD 0.00153f
C207 adder_4_1/adder_3_0/P2 GND 4.74e-20
C208 B12 VDD 0.0415f
C209 adder_4_1/CI adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 3.27e-22
C210 S4 S3 -9.65e-20
C211 adder_4_1/CI adder_4_2/adder_3_0/P2 4.97e-20
C212 adder_4_2/adder_3_0/P3 adder_4_3/adder_3_0/G3 2.38e-20
C213 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/P2 2.19e-20
C214 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S12 7.81e-20
C215 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 0.00903f
C216 adder_4_0/adder_3_0/P1 GND -1.14e-31
C217 adder_4_1/adder_3_0/P2 A11 1.97e-19
C218 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_0/adder_3_0/P2 5.27e-22
C219 adder_4_2/adder_2_0/G4 S7 2.25e-20
C220 B12 GND 0.00216f
C221 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# B16 1.9e-21
C222 adder_4_1/CI B6 5.55e-35
C223 adder_4_2/adder_2_0/G4 S6 1.98e-20
C224 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 2.53e-19
C225 adder_4_3/adder_3_0/G2 GND 1.6e-20
C226 adder_4_3/adder_3_0/P3 GND 1.01e-20
C227 A5 CI 3.01e-20
C228 adder_4_2/adder_3_0/G1 VDD 0.0748f
C229 adder_4_0/adder_3_0/P1 A6 1.27e-19
C230 S12 adder_4_3/adder_3_0/P4 2.69e-20
C231 A11 B12 1.11e-34
C232 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B12 5.68e-20
C233 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD 4.95e-20
C234 adder_4_2/adder_3_0/G1 GND 6.38e-21
C235 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A6 1.76e-20
C236 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 1.42e-19
C237 adder_4_1/adder_3_0/P3 adder_4_0/adder_3_0/P3 1.88e-19
C238 S7 A12 0.00571f
C239 adder_4_1/CI S2 0.0018f
C240 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.4e-20
C241 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.18e-19
C242 S6 A12 1.69e-19
C243 A16 adder_4_2/adder_3_0/G2 1.02e-19
C244 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.77e-20
C245 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.46e-19
C246 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 7.69e-21
C247 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/P3 2.36e-20
C248 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_2/adder_3_0/G3 6.86e-21
C249 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_4_2/CI 8.76e-20
C250 B5 adder_4_0/adder_3_0/G1 5.49e-20
C251 B6 CI 8.69e-19
C252 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A12 3.71e-19
C253 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.91e-21
C254 A16 S11 0.00571f
C255 B8 VDD 0.0415f
C256 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.39e-19
C257 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B VDD 1.37e-19
C258 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_2/adder_3_0/P2 5.27e-22
C259 S12 VDD 2.91e-19
C260 B8 GND 0.0477f
C261 A16 adder_4_2/CI 5.12e-19
C262 adder_4_2/CI adder_4_2/adder_3_0/P4 3.66e-20
C263 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.39e-20
C264 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD 2.78e-20
C265 B10 adder_4_1/adder_3_0/G2 6.51e-20
C266 adder_4_1/adder_3_0/G3 A12 1.06e-19
C267 S12 GND 6.99e-20
C268 S5 adder_4_2/CI 2.87e-19
C269 A16 B13 5.55e-35
C270 S2 adder_4_1/adder_3_0/P3 1.88e-20
C271 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/P3 2.47e-20
C272 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 0.00903f
C273 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.53e-19
C274 adder_4_2/adder_3_0/P2 adder_4_3/CI 6.08e-19
C275 adder_4_2/CI adder_4_1/adder_3_0/G2 1.47e-19
C276 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_0/adder_3_0/P3 3.3e-19
C277 S5 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.6e-21
C278 adder_4_0/adder_3_0/G2 B5 1.61e-19
C279 adder_4_0/adder_3_0/G1 A5 9.55e-19
C280 adder_4_1/CI adder_4_1/adder_2_0/G4 3.53e-20
C281 adder_4_1/adder_2_0/G4 adder_4_0/adder_3_0/P4 3.69e-21
C282 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_3/CI 2.04e-20
C283 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.76e-20
C284 B16 adder_4_3/CI 0.279f
C285 adder_4_2/CI adder_4_2/adder_3_0/P3 3.24e-20
C286 B11 VDD 0.0408f
C287 adder_4_2/adder_3_0/G1 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 8.69e-22
C288 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.66e-19
C289 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.75e-20
C290 adder_4_1/CI adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.34e-20
C291 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/CI 3.7e-20
C292 B11 GND 0.00112f
C293 adder_4_2/adder_3_0/G3 VDD 5.85e-20
C294 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B16 0.00191f
C295 B6 adder_4_0/adder_3_0/P2 1.84e-19
C296 B16 adder_4_3/adder_3_0/G1 -6.94e-36
C297 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_1/adder_3_0/P1 2.06e-19
C298 VDD adder_4_1/adder_3_0/P4 1.01e-19
C299 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A10 4.4e-20
C300 A7 VDD 0.0409f
C301 adder_4_2/adder_3_0/G3 GND 5.02e-20
C302 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 4.06e-20
C303 adder_4_0/adder_3_0/G1 B6 7.06e-20
C304 GND adder_4_1/adder_3_0/P4 0.0441f
C305 A7 GND 8.93e-19
C306 adder_4_2/adder_3_0/P3 B14 0.00256f
C307 adder_4_3/CI S9 2.87e-19
C308 adder_4_2/CI S7 7.11e-33
C309 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_1/adder_3_0/G1 8.69e-22
C310 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD 5.65e-20
C311 B8 S1 2.42e-19
C312 adder_4_2/CI S6 0.0018f
C313 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B VDD 0.00738f
C314 adder_4_2/adder_3_0/P3 B15 2.06e-19
C315 A9 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.68e-19
C316 S5 B12 2.42e-19
C317 B8 S4 5.46e-19
C318 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S7 2.47e-20
C319 GND adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.41e-20
C320 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.15e-20
C321 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S6 2.19e-20
C322 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/P3 2.47e-20
C323 adder_4_0/adder_3_0/P1 adder_4_1/adder_3_0/G2 5.87e-21
C324 adder_4_2/adder_3_0/P1 VDD 0.00153f
C325 A16 adder_4_2/adder_3_0/G1 1.1e-19
C326 B12 adder_4_1/adder_3_0/G2 1.21e-19
C327 adder_4_3/adder_2_0/G4 S9 1.75e-20
C328 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.9e-19
C329 A8 adder_4_0/adder_3_0/G3 1.06e-19
C330 B8 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.37e-21
C331 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/P1 4.66e-20
C332 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.29e-19
C333 A14 VDD 0.0431f
C334 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B16 5.68e-20
C335 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_3/CI 6.87e-20
C336 B10 adder_4_1/adder_3_0/G3 6.79e-20
C337 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.15e-20
C338 A14 GND 4.78e-19
C339 adder_4_0/adder_3_0/G2 B6 6.51e-20
C340 adder_4_3/adder_3_0/G2 adder_4_2/adder_3_0/P3 3.43e-21
C341 adder_4_3/adder_3_0/P3 adder_4_2/adder_3_0/P3 1.88e-19
C342 GND adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 1.01e-20
C343 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.68e-20
C344 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.01e-20
C345 A13 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.68e-19
C346 adder_4_1/adder_3_0/G3 adder_4_2/CI 1.54e-19
C347 adder_4_1/CI VDD 0.156f
C348 adder_4_0/adder_3_0/P4 VDD 1.01e-19
C349 B15 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.7e-20
C350 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 9.5e-20
C351 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# A12 3.19e-20
C352 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.43e-20
C353 B6 A5 1.11e-34
C354 A10 VDD 0.0431f
C355 adder_4_1/CI GND 0.101f
C356 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 9.5e-20
C357 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# GND 1.01e-20
C358 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/P1 1.07e-21
C359 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A12 3.19e-20
C360 A10 GND 4.78e-19
C361 S1 adder_4_1/adder_3_0/P4 1.83e-20
C362 adder_4_1/CI A11 2.75e-19
C363 B6 adder_4_0/adder_3_0/P3 0.00256f
C364 S1 A7 1.1e-19
C365 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.19e-22
C366 A12 B9 5.55e-35
C367 B12 S7 4.77e-19
C368 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_3/CI 3.7e-20
C369 B12 S6 3.18e-19
C370 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 7.91e-21
C371 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.91e-21
C372 S4 adder_4_1/adder_3_0/P4 2.69e-20
C373 B7 adder_4_0/adder_3_0/G3 9.04e-20
C374 A16 S12 3.33e-19
C375 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/P2 2.53e-19
C376 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.34e-20
C377 adder_4_3/CI adder_4_3/adder_3_0/P4 3.66e-20
C378 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.46e-19
C379 adder_4_2/adder_3_0/G2 A15 7.47e-20
C380 adder_4_2/adder_3_0/P2 B16 4.43e-19
C381 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.68e-20
C382 CI VDD 0.0691f
C383 adder_4_1/adder_3_0/G1 VDD 0.0748f
C384 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 3.19e-20
C385 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 0.00903f
C386 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 2.08e-19
C387 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.19e-22
C388 adder_4_1/adder_3_0/P3 VDD 0.00144f
C389 S8 A12 3.33e-19
C390 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A8 4.77e-20
C391 CI GND 3.79e-20
C392 adder_4_1/adder_3_0/G1 GND 6.38e-21
C393 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_1/adder_3_0/P1 5.99e-21
C394 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 7.69e-21
C395 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A15 6.15e-20
C396 adder_4_1/adder_3_0/P3 GND 1.01e-20
C397 A11 adder_4_1/adder_3_0/G1 8.1e-20
C398 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.32e-20
C399 CI A6 1.92e-19
C400 B8 adder_4_0/adder_2_0/G4 1.47e-21
C401 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 7.69e-21
C402 adder_4_1/adder_3_0/P1 B9 8.38e-20
C403 B12 adder_4_1/adder_3_0/G3 1.27e-19
C404 A15 adder_4_2/CI 2.75e-19
C405 A11 adder_4_1/adder_3_0/P3 2.29e-19
C406 B11 S5 8.93e-20
C407 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/P3 1.33e-20
C408 A16 adder_4_2/adder_3_0/G3 1.06e-19
C409 adder_4_1/CI S1 2.87e-19
C410 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# S9 5.99e-21
C411 B11 adder_4_1/adder_3_0/G2 8.67e-20
C412 S5 adder_4_2/adder_3_0/G3 1.85e-20
C413 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S10 1.18e-20
C414 B16 S9 2.42e-19
C415 adder_4_3/CI VDD 0.087f
C416 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.19e-20
C417 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.01e-20
C418 adder_4_1/CI adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.77e-21
C419 adder_4_3/CI GND 0.04f
C420 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_4_2/CI 2.04e-20
C421 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B7 4.06e-20
C422 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B VDD 0.00738f
C423 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_2/CI 4.64e-20
C424 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B14 2.01e-20
C425 adder_4_3/adder_3_0/G1 VDD 2.84e-32
C426 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_3/adder_3_0/G2 4.9e-21
C427 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S3 5.56e-20
C428 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.01e-20
C429 adder_4_0/adder_3_0/P2 VDD 9.04e-19
C430 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B15 2.7e-20
C431 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND 1.39e-20
C432 A16 adder_4_2/adder_3_0/P1 2.81e-19
C433 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B GND 3.41e-20
C434 B10 B9 -4.44e-34
C435 adder_4_3/adder_3_0/G1 GND 6.38e-21
C436 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00265f
C437 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A8 4.77e-20
C438 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 7.69e-21
C439 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B16 5.68e-20
C440 GND adder_4_0/adder_3_0/P2 -5.68e-32
C441 S10 B15 3.58e-19
C442 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 4.64e-20
C443 adder_4_3/adder_2_0/G4 GND 4.83e-20
C444 adder_4_0/adder_3_0/G1 VDD 0.0748f
C445 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.52e-21
C446 S1 adder_4_1/adder_3_0/P3 1.67e-20
C447 A6 adder_4_0/adder_3_0/P2 1.62e-19
C448 adder_4_0/adder_3_0/G1 GND 5.68e-32
C449 B11 S6 3.58e-19
C450 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# A12 3.39e-20
C451 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B VDD 1.37e-19
C452 A9 adder_4_1/adder_3_0/P1 2.83e-20
C453 B5 VDD 0.0449f
C454 A8 S3 0.00571f
C455 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# B16 8.75e-20
C456 adder_4_0/adder_3_0/G1 A6 6.2e-20
C457 S2 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 1.82e-19
C458 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.15e-20
C459 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.9e-20
C460 B5 GND 1.84e-19
C461 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD 5.51e-20
C462 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B VDD 0.00738f
C463 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.8e-21
C464 A15 adder_4_2/adder_3_0/G1 8.1e-20
C465 A14 adder_4_2/adder_3_0/P3 4.46e-20
C466 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.34e-20
C467 adder_4_3/adder_3_0/P3 S10 1.88e-20
C468 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.92e-22
C469 adder_4_1/CI adder_4_1/adder_3_0/G2 6.94e-36
C470 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 7.69e-21
C471 S2 adder_4_1/adder_2_0/G4 1.98e-20
C472 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B GND 3.41e-20
C473 adder_4_0/adder_3_0/G2 VDD 4.62e-20
C474 adder_4_1/CI adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.7e-20
C475 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B7 4.21e-20
C476 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S8 7.81e-20
C477 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.18e-20
C478 adder_4_1/adder_3_0/G2 A10 5.72e-20
C479 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-19
C480 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B12 3.81e-20
C481 B11 adder_4_1/adder_3_0/G3 9.04e-20
C482 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.75e-20
C483 A5 VDD 0.0675f
C484 B10 A9 1.11e-34
C485 B5 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.08e-21
C486 adder_4_0/adder_3_0/G2 A6 5.72e-20
C487 adder_4_1/CI adder_4_0/adder_2_0/G4 1.64e-21
C488 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.81e-20
C489 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S9 6.6e-21
C490 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 5e-21
C491 A5 GND 1.99e-19
C492 adder_4_1/adder_3_0/P1 A12 2.81e-19
C493 adder_4_0/adder_3_0/P3 VDD 0.00144f
C494 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.76e-20
C495 CI adder_4_1/adder_3_0/G2 8.7e-21
C496 S9 adder_4_3/adder_3_0/P4 1.83e-20
C497 GND adder_4_0/adder_3_0/P3 1.14e-31
C498 adder_4_2/adder_3_0/P2 VDD 9.04e-19
C499 adder_4_1/adder_3_0/G3 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.18e-20
C500 A6 adder_4_0/adder_3_0/P3 4.46e-20
C501 adder_4_2/adder_3_0/P2 GND 4.74e-20
C502 B6 VDD 0.0407f
C503 B12 S8 5.46e-19
C504 B16 VDD 0.0415f
C505 adder_4_2/CI adder_4_2/adder_2_0/G4 3.53e-20
C506 adder_4_0/adder_3_0/P1 A8 2.81e-19
C507 adder_4_2/adder_3_0/P3 adder_4_1/adder_3_0/P3 1.88e-19
C508 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.32e-20
C509 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# GND 1.66e-20
C510 B6 GND 6.79e-19
C511 A5 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.22e-19
C512 A16 adder_4_3/CI 0.00128f
C513 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S3 2.47e-20
C514 B16 GND 0.00216f
C515 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A8 3.19e-20
C516 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/P3 3.44e-19
C517 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_3/adder_3_0/G3 6.86e-21
C518 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.42e-19
C519 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0011f
C520 S2 VDD 3.45e-19
C521 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.46e-19
C522 A16 adder_4_3/adder_3_0/G1 -1.39e-35
C523 adder_4_1/CI adder_4_1/adder_3_0/G3 9.03e-20
C524 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/P2 2.08e-20
C525 adder_4_2/CI A12 0.00128f
C526 S2 GND 0.0389f
C527 A15 adder_4_2/adder_3_0/G3 7.8e-20
C528 adder_4_3/adder_2_0/G4 adder_4_2/adder_3_0/P4 3.69e-21
C529 S9 VDD 8.75e-19
C530 adder_4_1/adder_3_0/G3 A10 8.92e-19
C531 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_2/adder_3_0/G3 2.84e-32
C532 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C533 adder_4_3/CI adder_4_2/adder_3_0/P3 7.78e-19
C534 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.78e-20
C535 adder_4_2/adder_3_0/G2 adder_4_1/adder_3_0/P1 5.87e-21
C536 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/P2 6.64e-21
C537 adder_4_3/CI adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.77e-21
C538 adder_4_0/adder_3_0/P1 B7 2.28e-19
C539 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.7e-20
C540 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B7 2.7e-20
C541 B10 adder_4_1/adder_3_0/P1 1.48e-19
C542 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.01e-20
C543 CI adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 9.5e-20
C544 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 5.65e-20
C545 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.71e-19
C546 A15 adder_4_2/adder_3_0/P1 1.89e-19
C547 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.7e-20
C548 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.4e-20
C549 adder_4_2/CI adder_4_1/adder_3_0/P1 4.71e-19
C550 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_4_2/CI 3.27e-22
C551 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# VDD 4.75e-20
C552 B8 adder_4_0/adder_3_0/G3 1.27e-19
C553 adder_4_3/CI adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 4.64e-20
C554 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.9e-19
C555 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.19e-20
C556 adder_4_1/adder_3_0/P2 A12 3.39e-19
C557 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# S3 1.39e-20
C558 adder_4_1/adder_2_0/G4 GND 6.02e-20
C559 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.19e-22
C560 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 6.83e-22
C561 adder_4_2/adder_3_0/G2 adder_4_2/CI 6.94e-36
C562 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.8e-20
C563 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B VDD 0.0303f
C564 adder_4_2/adder_3_0/P3 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.97e-20
C565 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.14e-19
C566 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.27e-22
C567 S2 S4 -9.65e-20
C568 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# GND 1.39e-20
C569 adder_4_2/adder_3_0/G2 B13 1.61e-19
C570 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/P3 2.47e-20
C571 adder_4_2/adder_3_0/G1 A12 -1.39e-35
C572 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.52e-21
C573 B8 B7 2.22e-34
C574 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S8 1.16e-19
C575 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# S10 1.82e-19
C576 B10 adder_4_2/CI 5.55e-35
C577 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.15e-20
C578 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.9e-21
C579 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 3.96e-19
C580 S11 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.56e-20
C581 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A12 4.77e-20
C582 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.72e-21
C583 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.28e-21
C584 adder_4_3/adder_3_0/P4 GND 4.46e-20
C585 A16 adder_4_2/adder_3_0/P2 3.39e-19
C586 adder_4_2/adder_3_0/G2 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.9e-21
C587 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B B14 2.79e-20
C588 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/P3 3.43e-21
C589 adder_4_2/adder_3_0/G2 B14 6.51e-20
C590 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B13 4.08e-21
C591 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B B15 2.72e-21
C592 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.7e-20
C593 adder_4_2/adder_3_0/G2 B15 8.67e-20
C594 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B15 4.21e-20
C595 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/P3 3.44e-19
C596 adder_4_1/adder_3_0/G3 adder_4_0/adder_3_0/P2 4e-21
C597 B12 adder_4_1/adder_3_0/P1 3.59e-19
C598 B16 adder_4_2/adder_3_0/P4 1.24e-19
C599 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.52e-20
C600 A7 adder_4_0/adder_3_0/G3 7.8e-20
C601 adder_4_2/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.7e-20
C602 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# A10 3.9e-19
C603 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.19e-20
C604 adder_4_2/CI B13 1.09e-19
C605 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# B12 2.93e-22
C606 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 6.83e-22
C607 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0011f
C608 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_4_3/CI 6.93e-21
C609 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B14 5.78e-20
C610 adder_4_1/CI B9 1.09e-19
C611 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.68e-20
C612 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A13 1.22e-19
C613 adder_4_2/adder_3_0/G2 adder_4_1/adder_3_0/P2 6.64e-21
C614 adder_4_1/CI adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 2.04e-20
C615 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_0/adder_3_0/G3 2.84e-32
C616 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B15 1.18e-19
C617 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.76e-20
C618 adder_4_2/adder_3_0/G1 adder_4_1/adder_3_0/P1 7.91e-22
C619 adder_4_2/CI B14 8.69e-19
C620 S1 adder_4_1/adder_2_0/G4 1.75e-20
C621 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_3/adder_3_0/G1 8.69e-22
C622 A13 adder_4_2/CI 3.01e-20
C623 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 7.91e-21
C624 adder_4_2/CI B15 3.65e-19
C625 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/P3 1.33e-20
C626 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.52e-20
C627 adder_4_3/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.7e-20
C628 A16 S9 1.3e-19
C629 B16 adder_4_2/adder_3_0/P3 5.72e-19
C630 S12 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 1.16e-19
C631 adder_4_1/adder_3_0/P2 B10 1.84e-19
C632 GND VDD 0.385f
C633 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/CI 5.01e-20
C634 B16 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.37e-21
C635 adder_4_3/adder_3_0/P1 adder_4_2/CI 2.44e-20
C636 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.52e-21
C637 adder_4_1/adder_3_0/P2 adder_4_2/CI 9.44e-19
C638 adder_4_1/CI A8 0.00128f
C639 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S2 5.48e-20
C640 A15 adder_4_3/CI 0.00338f
C641 A11 VDD 0.0409f
C642 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 5.65e-20
C643 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# GND 1.39e-20
C644 A6 VDD 0.0431f
C645 adder_4_2/adder_2_0/G4 adder_4_1/adder_3_0/P4 3.69e-21
C646 adder_4_3/CI adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.64e-20
C647 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S4 1.16e-19
C648 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.7e-20
C649 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00977f
C650 A13 B14 1.11e-34
C651 adder_4_1/adder_3_0/G1 B9 5.49e-20
C652 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C653 B12 adder_4_2/CI 0.279f
C654 B9 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.56e-20
C655 A11 GND 8.93e-19
C656 A6 GND 4.78e-19
C657 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S8 2.71e-19
C658 adder_4_1/CI adder_4_0/adder_3_0/G3 1.54e-19
C659 B1 VDD 5.67e-22
C660 adder_4_3/adder_3_0/G2 adder_4_2/CI 8.7e-21
C661 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.39e-20
C662 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-19
C663 adder_4_3/CI S10 0.0018f
C664 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# GND 1.66e-20
C665 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 4.77e-20
C666 adder_4_0/adder_3_0/P1 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 5.99e-21
C667 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A11 3.5e-20
C668 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.92e-22
C669 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.2e-20
C670 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.81e-20
C671 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B VDD 0.0303f
C672 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A7 3.5e-20
C673 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.68e-20
C674 adder_4_1/adder_3_0/G3 adder_4_0/adder_3_0/P3 2.38e-20
C675 adder_4_3/adder_3_0/P2 GND 4.74e-20
C676 adder_4_3/adder_2_0/G4 S10 1.98e-20
C677 adder_4_1/CI A9 3.01e-20
C678 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.44e-19
C679 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.39e-35
C680 adder_4_2/adder_3_0/G1 B13 5.49e-20
C681 CI A8 5.12e-19
C682 A8 adder_4_1/adder_3_0/G1 -1.39e-35
C683 adder_4_1/CI B7 7.44e-19
C684 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.4e-20
C685 adder_4_3/adder_3_0/G2 B15 1.39e-35
C686 B8 S3 4.77e-19
C687 adder_4_2/adder_3_0/G1 B14 7.06e-20
C688 S1 VDD 8.75e-19
C689 B11 adder_4_1/adder_3_0/P1 2.28e-19
C690 adder_4_2/adder_3_0/G1 A13 9.55e-19
C691 adder_4_0/adder_3_0/P1 adder_4_1/adder_3_0/P2 1.07e-21
C692 adder_4_2/adder_3_0/G1 B15 9.39e-20
C693 adder_4_1/adder_3_0/P2 B12 4.43e-19
C694 S4 VDD 2.91e-19
C695 S1 GND 0.036f
C696 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C697 S4 GND 0.071f
C698 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_2/CI 3.96e-19
C699 adder_4_1/adder_3_0/G1 A9 9.55e-19
C700 A9 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.25e-19
C701 B11 adder_4_2/adder_3_0/G2 1.39e-35
C702 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.87e-20
C703 adder_4_1/CI A12 5.12e-19
C704 adder_4_1/CI adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.7e-20
C705 CI B7 3.65e-19
C706 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# B16 2.93e-22
C707 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# B12 8.75e-20
C708 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A7 2.46e-19
C709 adder_4_2/adder_3_0/G1 B12 -6.94e-36
C710 adder_4_1/adder_3_0/P1 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.81e-20
C711 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.75e-20
C712 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD 5.51e-20
C713 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.68e-20
C714 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.22e-19
C715 B11 B10 4.44e-34
C716 A8 adder_4_0/adder_3_0/P2 3.39e-19
C717 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B13 1.56e-20
C718 S3 adder_4_1/adder_3_0/P4 2.35e-20
C719 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B9 0.00399f
C720 A15 adder_4_2/adder_3_0/P2 1.97e-19
C721 B11 adder_4_2/CI 7.44e-19
C722 adder_4_0/adder_3_0/G1 A8 1.1e-19
C723 A16 VDD 0.0408f
C724 adder_4_2/adder_3_0/P4 VDD 1.01e-19
C725 adder_4_2/CI adder_4_2/adder_3_0/G3 4.85e-20
C726 S5 VDD 8.75e-19
C727 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_3/CI 3.96e-19
C728 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B14 2.01e-20
C729 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# GND 8.39e-19
C730 A15 B16 1.11e-34
C731 A13 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.25e-19
C732 A16 GND 0.00154f
C733 adder_4_2/adder_3_0/P4 GND 4.46e-20
C734 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B15 2.7e-20
C735 adder_4_1/adder_3_0/G1 A12 1.1e-19
C736 B8 adder_4_0/adder_3_0/P1 3.59e-19
C737 A12 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 3.19e-20
C738 adder_4_1/CI adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 2.04e-20
C739 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_2/adder_3_0/P1 6.6e-21
C740 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.81e-20
C741 B5 A8 5.55e-35
C742 adder_4_1/adder_3_0/G2 VDD 4.62e-20
C743 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.53e-19
C744 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_1/adder_3_0/P1 6.6e-21
C745 adder_4_1/adder_3_0/P3 A12 4.13e-19
C746 A14 adder_4_2/adder_3_0/G2 5.72e-20
C747 B16 S10 3.18e-19
C748 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B8 3.81e-20
C749 S1 S4 -9.65e-20
C750 A10 adder_4_1/adder_3_0/P1 1.27e-19
C751 S5 A11 1.1e-19
C752 adder_4_1/adder_3_0/G2 GND 1.6e-20
C753 S9 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.6e-21
C754 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.44e-19
C755 S5 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 5.99e-21
C756 adder_4_3/CI adder_4_2/adder_2_0/G4 1.64e-21
C757 adder_4_2/adder_3_0/P3 VDD 0.00144f
C758 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_3/CI 1.39e-35
C759 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# GND 1.17e-20
C760 B7 adder_4_0/adder_3_0/P2 3.03e-19
C761 A11 adder_4_1/adder_3_0/G2 7.47e-20
C762 adder_4_2/adder_3_0/G3 B14 6.79e-20
C763 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 7.69e-21
C764 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.22e-19
C765 adder_4_1/CI adder_4_2/adder_3_0/G2 8.7e-21
C766 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.4e-20
C767 adder_4_2/adder_3_0/P3 GND 1.01e-20
C768 adder_4_0/adder_3_0/G2 A8 1.02e-19
C769 adder_4_2/adder_3_0/G3 B15 9.04e-20
C770 A15 S9 1.1e-19
C771 adder_4_2/CI adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.77e-21
C772 adder_4_0/adder_3_0/G1 B7 9.39e-20
C773 B11 adder_4_1/adder_3_0/P2 3.03e-19
C774 A14 adder_4_2/CI 1.92e-19
C775 adder_4_1/CI S3 7.11e-33
C776 A2 VDD 1.54e-22
C777 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# GND 1.17e-20
C778 adder_4_3/adder_2_0/G4 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.82e-21
C779 B13 adder_4_2/adder_3_0/P1 8.38e-20
C780 CI adder_4_1/adder_3_0/P1 2.44e-20
C781 adder_4_3/CI adder_4_3/adder_3_0/G3 4.85e-20
C782 adder_4_1/CI B10 8.69e-19
C783 adder_4_1/adder_3_0/P2 adder_4_2/adder_3_0/G3 4e-21
C784 A9 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.79e-20
C785 S7 VDD 2.72e-19
C786 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# S7 1.39e-20
C787 S6 VDD 3.45e-19
C788 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_3_0/G3 3.18e-20
C789 A8 adder_4_0/adder_3_0/P3 4.13e-19
C790 adder_4_1/CI adder_4_2/CI 0.0496f
C791 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.5e-20
C792 CI adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# 8.76e-20
C793 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/P3 2.36e-20
C794 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD 2.78e-20
C795 adder_4_2/adder_3_0/P1 B14 1.48e-19
C796 adder_4_2/adder_2_0/G4 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 9.08e-21
C797 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_4_2/CI 2.13e-21
C798 A13 adder_4_2/adder_3_0/P1 2.83e-20
C799 GND S6 3.33e-22
C800 adder_4_0/adder_3_0/P1 A7 1.89e-19
C801 B12 adder_4_1/adder_3_0/P4 1.24e-19
C802 B15 adder_4_2/adder_3_0/P1 2.28e-19
C803 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD 5.51e-20
C804 adder_4_1/adder_3_0/P2 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.15e-20
C805 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S4 2.71e-19
C806 B8 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.9e-21
C807 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.74e-19
C808 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/adder_3_0/P1 5.99e-21
C809 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_4_3/CI 4.91e-21
C810 A11 S6 3.71e-20
C811 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.21e-20
C812 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A7 2.32e-20
C813 S2 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 1.18e-20
C814 adder_4_2/adder_3_0/G2 adder_4_1/adder_3_0/P3 3.43e-21
C815 adder_4_0/adder_3_0/G2 B7 8.67e-20
C816 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/P1 4.66e-20
C817 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.81e-20
C818 adder_4_1/adder_3_0/P2 adder_4_2/adder_3_0/P1 0.00296f
C819 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S1 6.6e-21
C820 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B A12 1.4e-20
C821 B10 adder_4_1/adder_3_0/G1 7.06e-20
C822 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.01e-20
C823 B6 adder_4_0/adder_3_0/G3 6.79e-20
C824 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# 8.76e-20
C825 adder_4_1/adder_3_0/G3 VDD 5.85e-20
C826 B10 adder_4_1/adder_3_0/P3 0.00256f
C827 B12 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.37e-21
C828 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# GND 1.39e-20
C829 adder_4_3/adder_3_0/G2 adder_4_2/adder_3_0/P1 5.87e-21
C830 adder_4_2/CI adder_4_1/adder_3_0/G1 1.58e-19
C831 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 4.64e-20
C832 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_2/adder_3_0/P3 3.3e-19
C833 adder_4_1/adder_3_0/G3 GND 5.02e-20
C834 adder_4_0/adder_3_0/P1 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.6e-21
C835 B7 adder_4_0/adder_3_0/P3 2.06e-19
C836 adder_4_2/CI adder_4_1/adder_3_0/P3 7.78e-19
C837 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A12 0.0011f
C838 S2 A8 1.69e-19
C839 adder_4_1/adder_3_0/P1 adder_4_0/adder_3_0/P2 0.00296f
C840 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/P2 2.53e-19
C841 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# GND 1.39e-20
C842 CI adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.52e-20
C843 adder_4_0/adder_3_0/P1 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.06e-19
C844 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S10 2.19e-20
C845 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/CI 5.9e-20
C846 A11 adder_4_1/adder_3_0/G3 7.8e-20
C847 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# S6 1.82e-19
C848 adder_4_2/adder_3_0/G2 adder_4_3/CI 1.47e-19
C849 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.8e-21
C850 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_3/CI 7.44e-19
C851 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.6e-19
C852 adder_4_1/CI adder_4_0/adder_3_0/P1 4.71e-19
C853 A14 adder_4_2/adder_3_0/G1 6.2e-20
C854 adder_4_1/adder_3_0/P2 A10 1.62e-19
C855 adder_4_3/adder_3_0/P4 S10 2.06e-20
C856 adder_4_1/CI B12 7.74e-19
C857 B8 A7 1.11e-34
C858 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# B12 1.9e-21
C859 adder_4_1/adder_3_0/P3 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.3e-19
C860 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 9.13e-20
C861 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 4.64e-20
C862 adder_4_3/CI S11 7.11e-33
C863 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.34e-20
C864 adder_4_3/adder_2_0/G4 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 9.08e-21
C865 S5 adder_4_2/adder_3_0/P4 1.83e-20
C866 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_3/CI 2.56e-19
C867 S12 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 2.71e-19
C868 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND 1.39e-20
C869 adder_4_1/adder_3_0/G3 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.86e-21
C870 adder_4_1/CI adder_4_2/adder_3_0/G1 0.0031f
C871 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.81e-20
C872 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00191f
C873 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.32e-20
C874 adder_4_2/CI adder_4_3/CI 0.0496f
C875 B16 adder_4_2/adder_2_0/G4 1.47e-21
C876 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD -5.68e-32
C877 adder_4_3/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 2.04e-20
C878 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# B16 2.14e-19
C879 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B9 4.08e-21
C880 adder_4_3/adder_2_0/G4 S11 2.25e-20
C881 adder_4_1/adder_3_0/P2 CI 4.97e-20
C882 S2 B7 3.58e-19
C883 A16 adder_4_2/adder_3_0/P3 4.13e-19
C884 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# GND 1.17e-20
C885 adder_4_2/adder_3_0/P2 adder_4_3/adder_3_0/G3 4e-21
C886 adder_4_2/CI adder_4_3/adder_3_0/G1 0.0031f
C887 A15 VDD 0.0409f
C888 adder_4_0/adder_3_0/P1 adder_4_1/adder_3_0/G1 7.91e-22
C889 S5 adder_4_2/adder_3_0/P3 1.67e-20
C890 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 3.81e-20
C891 B12 adder_4_1/adder_3_0/G1 1.31e-19
C892 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B6 2.06e-22
C893 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD 5.65e-20
C894 S1 adder_4_1/adder_3_0/G3 1.85e-20
C895 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B13 0.00399f
C896 A15 GND 8.93e-19
C897 B12 adder_4_1/adder_3_0/P3 5.72e-19
C898 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/P2 1.18e-20
C899 S10 VDD 3.45e-19
C900 S5 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.6e-21
C901 adder_4_3/CI B14 5.55e-35
C902 adder_4_2/adder_3_0/G2 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00265f
C903 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.79e-20
C904 adder_4_3/CI B15 7.76e-19
C905 adder_4_1/CI B8 0.279f
C906 B8 adder_4_0/adder_3_0/P4 1.24e-19
C907 S10 GND 3.33e-22
C908 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.9e-20
C909 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B14 4.05e-19
C910 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.9e-20
C911 A13 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.79e-20
C912 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.76e-20
C913 adder_4_2/adder_3_0/P4 S7 2.35e-20
C914 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/P3 1.33e-20
C915 adder_4_1/CI adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 2.13e-21
C916 adder_4_2/adder_3_0/P4 S6 2.06e-20
C917 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B15 0.00977f
C918 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.05e-19
C919 S2 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.19e-20
C920 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.19e-20
C921 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD 5.65e-20
C922 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.22e-19
C923 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X B16 4.4e-21
C924 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 7.91e-21
C925 adder_4_1/CI adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 4.64e-20
C926 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# GND 1.76e-20
C927 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.32e-20
C928 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/P1 1.07e-21
C929 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-19
C930 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 3.2e-20
C931 S9 adder_4_3/adder_3_0/G3 1.85e-20
C932 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.433f
C933 adder_4_1/adder_2_0/G4 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.82e-21
C934 adder_4_3/adder_3_0/P1 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.81e-20
C935 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD 2.78e-20
C936 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# GND 1.39e-20
C937 adder_4_3/adder_3_0/G2 adder_4_3/CI 6.94e-36
C938 B9 VDD 0.0449f
C939 adder_4_3/adder_3_0/P3 adder_4_3/CI 3.24e-20
C940 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# A11 2.32e-20
C941 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A9 1.22e-19
C942 adder_4_1/adder_3_0/P2 adder_4_0/adder_3_0/P2 2.08e-20
C943 A14 adder_4_2/adder_3_0/G3 8.92e-19
C944 adder_4_0/adder_3_0/P1 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.66e-20
C945 adder_4_2/adder_3_0/P3 S6 1.88e-20
C946 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_2/adder_2_0/G4 3.82e-21
C947 GND B9 1.84e-19
C948 B8 CI 7.74e-19
C949 B8 adder_4_1/adder_3_0/G1 -6.94e-36
C950 adder_4_3/adder_3_0/G2 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00265f
C951 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 5e-21
C952 B11 adder_4_1/CI 3.65e-19
C953 adder_4_2/adder_3_0/G1 adder_4_3/CI 1.58e-19
C954 adder_4_3/adder_3_0/P3 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.97e-20
C955 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# GND 1.76e-20
C956 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.32e-20
C957 adder_4_2/adder_3_0/P2 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.6e-19
C958 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S6 5.48e-20
C959 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.92e-22
C960 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B15 2.9e-20
C961 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B B16 3.74e-19
C962 adder_4_2/adder_3_0/G2 B16 1.21e-19
C963 adder_4_1/CI adder_4_1/adder_3_0/P4 3.66e-20
C964 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B16 5.68e-20
C965 S8 VDD 2.91e-19
C966 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 9.13e-20
C967 adder_4_1/CI A7 0.00338f
C968 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C969 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C970 A2 0 0.553f
C971 B2 0 0.632f
C972 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C973 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C974 A1 0 0.469f
C975 B1 0 0.496f
C976 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C977 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C978 B4 0 1.05f
C979 A4 0 0.714f
C980 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C981 B3 0 0.683f
C982 A3 0 0.729f
C983 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C984 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C985 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C986 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C987 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C988 S3 0 0.226f
C989 adder_4_0/adder_3_0/P3 0 1.49f
C990 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C991 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C992 S2 0 0.212f
C993 adder_4_0/adder_3_0/P2 0 1.26f
C994 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C995 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C996 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C997 S1 0 0.285f
C998 adder_4_0/adder_3_0/P1 0 1.11f
C999 CI 0 2.13f
C1000 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1001 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1002 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1003 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1004 adder_4_0/adder_3_0/G3 0 0.718f
C1005 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1006 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1007 adder_4_0/adder_3_0/G2 0 0.642f
C1008 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1009 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1010 adder_4_0/adder_3_0/G1 0 0.527f
C1011 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1012 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1013 S4 0 0.305f
C1014 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1015 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1016 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1017 adder_4_0/adder_3_0/P4 0 1.62f
C1018 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1019 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1020 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1021 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1022 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1023 adder_4_0/adder_2_0/G4 0 0.596f
C1024 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1025 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1026 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1027 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1028 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1029 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1030 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1031 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1032 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1033 A14 0 0.547f
C1034 B14 0 0.627f
C1035 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1036 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1037 A13 0 0.45f
C1038 B13 0 0.484f
C1039 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1040 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1041 B16 0 1.05f
C1042 A16 0 0.714f
C1043 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C1044 B15 0 0.683f
C1045 A15 0 0.729f
C1046 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C1047 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C1048 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C1049 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1050 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1051 S15 0 0.233f
C1052 adder_4_3/adder_3_0/P3 0 1.49f
C1053 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1054 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1055 S14 0 0.212f
C1056 adder_4_3/adder_3_0/P2 0 1.26f
C1057 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C1058 VDD 0 71.6f
C1059 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1060 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1061 S13 0 0.285f
C1062 adder_4_3/adder_3_0/P1 0 1.11f
C1063 adder_4_3/CI 0 2.22f
C1064 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1065 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1066 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1067 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1068 adder_4_3/adder_3_0/G3 0 0.718f
C1069 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1070 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1071 adder_4_3/adder_3_0/G2 0 0.642f
C1072 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1073 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1074 adder_4_3/adder_3_0/G1 0 0.527f
C1075 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1076 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1077 S16 0 0.335f
C1078 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1079 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1080 adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1081 adder_4_3/adder_3_0/P4 0 1.62f
C1082 adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1083 CO 0 0.959f
C1084 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1085 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1086 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1087 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1088 adder_4_3/adder_2_0/G4 0 0.596f
C1089 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1090 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1091 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1092 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1093 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1094 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1095 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1096 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1097 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1098 A10 0 0.547f
C1099 B10 0 0.627f
C1100 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1101 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1102 A9 0 0.45f
C1103 B9 0 0.484f
C1104 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1105 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1106 B12 0 1.05f
C1107 A12 0 0.714f
C1108 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C1109 B11 0 0.683f
C1110 A11 0 0.729f
C1111 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C1112 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C1113 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C1114 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1115 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1116 S11 0 0.226f
C1117 adder_4_2/adder_3_0/P3 0 1.49f
C1118 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1119 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1120 S10 0 0.212f
C1121 adder_4_2/adder_3_0/P2 0 1.26f
C1122 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C1123 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1124 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1125 S9 0 0.285f
C1126 adder_4_2/adder_3_0/P1 0 1.11f
C1127 adder_4_2/CI 0 2.23f
C1128 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1129 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1130 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1131 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1132 adder_4_2/adder_3_0/G3 0 0.718f
C1133 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1134 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1135 adder_4_2/adder_3_0/G2 0 0.642f
C1136 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1137 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1138 adder_4_2/adder_3_0/G1 0 0.527f
C1139 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1140 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1141 S12 0 0.334f
C1142 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1143 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1144 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1145 adder_4_2/adder_3_0/P4 0 1.62f
C1146 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1147 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1148 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1149 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1150 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1151 adder_4_2/adder_2_0/G4 0 0.596f
C1152 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1153 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1154 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1155 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1156 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1157 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1158 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1159 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1160 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1161 A6 0 0.547f
C1162 B6 0 0.627f
C1163 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1164 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1165 A5 0 0.45f
C1166 B5 0 0.484f
C1167 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1168 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1169 B8 0 1.05f
C1170 A8 0 0.714f
C1171 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C1172 B7 0 0.683f
C1173 A7 0 0.729f
C1174 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C1175 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C1176 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C1177 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1178 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1179 S7 0 0.226f
C1180 adder_4_1/adder_3_0/P3 0 1.49f
C1181 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1182 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1183 GND 0 34.5f
C1184 S6 0 0.212f
C1185 adder_4_1/adder_3_0/P2 0 1.26f
C1186 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C1187 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1188 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1189 S5 0 0.285f
C1190 adder_4_1/adder_3_0/P1 0 1.11f
C1191 adder_4_1/CI 0 2.22f
C1192 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1193 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1194 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1195 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1196 adder_4_1/adder_3_0/G3 0 0.718f
C1197 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1198 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1199 adder_4_1/adder_3_0/G2 0 0.642f
C1200 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1201 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1202 adder_4_1/adder_3_0/G1 0 0.527f
C1203 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1204 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1205 S8 0 0.334f
C1206 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1207 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1208 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1209 adder_4_1/adder_3_0/P4 0 1.62f
C1210 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1211 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1212 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1213 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1214 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1215 adder_4_1/adder_2_0/G4 0 0.596f
C1216 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1217 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1218 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1219 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1220 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1221 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1222 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

